--------------------------------------------------------------------------------
--                          Compressor_6_3_F800_uid6
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_F800_uid6 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_F800_uid6 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_14_3_F800_uid10
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_F800_uid10 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_F800_uid10 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_3_2_F800_uid16
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_F800_uid16 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_F800_uid16 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_5_3_F800_uid98
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_F800_uid98 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_F800_uid98 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_23_3_F800_uid136
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_F800_uid136 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_F800_uid136 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_21_F800_uid186
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_21_F800_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(20 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntAdder_21_F800_uid186 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3 :  std_logic;
signal X_1, X_1_d1 :  std_logic_vector(15 downto 0);
signal Y_1, Y_1_d1 :  std_logic_vector(15 downto 0);
signal S_1 :  std_logic_vector(15 downto 0);
signal R_1, R_1_d1 :  std_logic_vector(14 downto 0);
signal Cin_2, Cin_2_d1 :  std_logic;
signal X_2, X_2_d1, X_2_d2 :  std_logic_vector(6 downto 0);
signal Y_2, Y_2_d1, Y_2_d2 :  std_logic_vector(6 downto 0);
signal S_2 :  std_logic_vector(6 downto 0);
signal R_2 :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
            R_1_d1 <=  R_1;
            Cin_2_d1 <=  Cin_2;
            X_2_d1 <=  X_2;
            X_2_d2 <=  X_2_d1;
            Y_2_d1 <=  Y_2;
            Y_2_d2 <=  Y_2_d1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(14 downto 0);
   Y_1 <= '0' & Y(14 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d3;
   R_1 <= S_1(14 downto 0);
   Cin_2 <= S_1(15);
   X_2 <= '0' & X(20 downto 15);
   Y_2 <= '0' & Y(20 downto 15);
   S_2 <= X_2_d2 + Y_2_d2 + Cin_2_d1;
   R_2 <= S_2(5 downto 0);
   R <= R_2 & R_1_d1 ;
end architecture;

--------------------------------------------------------------------------------
--                       IntMultiAdder_U20_10_F800_uid2
-- VHDL generated for Virtex6 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0 X1 X2 X3 X4 X5 X6 X7 X8 X9
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiAdder_U20_10_F800_uid2 is
    port (clk : in std_logic;
          R : out  std_logic_vector(23 downto 0);
          X0 : in  std_logic_vector(19 downto 0);
          X1 : in  std_logic_vector(19 downto 0);
          X2 : in  std_logic_vector(19 downto 0);
          X3 : in  std_logic_vector(19 downto 0);
          X4 : in  std_logic_vector(19 downto 0);
          X5 : in  std_logic_vector(19 downto 0);
          X6 : in  std_logic_vector(19 downto 0);
          X7 : in  std_logic_vector(19 downto 0);
          X8 : in  std_logic_vector(19 downto 0);
          X9 : in  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of IntMultiAdder_U20_10_F800_uid2 is
   component Compressor_6_3_F800_uid6 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_F800_uid10 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_F800_uid16 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_5_3_F800_uid98 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_23_3_F800_uid136 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_21_F800_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(20 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(20 downto 0)   );
   end component;

signal iX0 :  unsigned(19-0 downto 0);
signal bh3_w0_0 :  std_logic;
signal bh3_w1_0 :  std_logic;
signal bh3_w2_0 :  std_logic;
signal bh3_w3_0 :  std_logic;
signal bh3_w4_0 :  std_logic;
signal bh3_w5_0 :  std_logic;
signal bh3_w6_0 :  std_logic;
signal bh3_w7_0 :  std_logic;
signal bh3_w8_0 :  std_logic;
signal bh3_w9_0 :  std_logic;
signal bh3_w10_0 :  std_logic;
signal bh3_w11_0 :  std_logic;
signal bh3_w12_0 :  std_logic;
signal bh3_w13_0 :  std_logic;
signal bh3_w14_0 :  std_logic;
signal bh3_w15_0 :  std_logic;
signal bh3_w16_0 :  std_logic;
signal bh3_w17_0 :  std_logic;
signal bh3_w18_0 :  std_logic;
signal bh3_w19_0 :  std_logic;
signal iX1 :  unsigned(19-0 downto 0);
signal bh3_w0_1 :  std_logic;
signal bh3_w1_1 :  std_logic;
signal bh3_w2_1 :  std_logic;
signal bh3_w3_1 :  std_logic;
signal bh3_w4_1 :  std_logic;
signal bh3_w5_1 :  std_logic;
signal bh3_w6_1 :  std_logic;
signal bh3_w7_1 :  std_logic;
signal bh3_w8_1 :  std_logic;
signal bh3_w9_1 :  std_logic;
signal bh3_w10_1 :  std_logic;
signal bh3_w11_1 :  std_logic;
signal bh3_w12_1 :  std_logic;
signal bh3_w13_1 :  std_logic;
signal bh3_w14_1 :  std_logic;
signal bh3_w15_1 :  std_logic;
signal bh3_w16_1 :  std_logic;
signal bh3_w17_1 :  std_logic;
signal bh3_w18_1 :  std_logic;
signal bh3_w19_1 :  std_logic;
signal iX2 :  unsigned(19-0 downto 0);
signal bh3_w0_2 :  std_logic;
signal bh3_w1_2 :  std_logic;
signal bh3_w2_2 :  std_logic;
signal bh3_w3_2 :  std_logic;
signal bh3_w4_2 :  std_logic;
signal bh3_w5_2 :  std_logic;
signal bh3_w6_2 :  std_logic;
signal bh3_w7_2 :  std_logic;
signal bh3_w8_2 :  std_logic;
signal bh3_w9_2 :  std_logic;
signal bh3_w10_2 :  std_logic;
signal bh3_w11_2 :  std_logic;
signal bh3_w12_2 :  std_logic;
signal bh3_w13_2 :  std_logic;
signal bh3_w14_2 :  std_logic;
signal bh3_w15_2 :  std_logic;
signal bh3_w16_2 :  std_logic;
signal bh3_w17_2 :  std_logic;
signal bh3_w18_2 :  std_logic;
signal bh3_w19_2 :  std_logic;
signal iX3 :  unsigned(19-0 downto 0);
signal bh3_w0_3 :  std_logic;
signal bh3_w1_3 :  std_logic;
signal bh3_w2_3 :  std_logic;
signal bh3_w3_3 :  std_logic;
signal bh3_w4_3 :  std_logic;
signal bh3_w5_3 :  std_logic;
signal bh3_w6_3 :  std_logic;
signal bh3_w7_3 :  std_logic;
signal bh3_w8_3 :  std_logic;
signal bh3_w9_3 :  std_logic;
signal bh3_w10_3 :  std_logic;
signal bh3_w11_3 :  std_logic;
signal bh3_w12_3 :  std_logic;
signal bh3_w13_3 :  std_logic;
signal bh3_w14_3 :  std_logic;
signal bh3_w15_3 :  std_logic;
signal bh3_w16_3 :  std_logic;
signal bh3_w17_3 :  std_logic;
signal bh3_w18_3 :  std_logic;
signal bh3_w19_3 :  std_logic;
signal iX4 :  unsigned(19-0 downto 0);
signal bh3_w0_4 :  std_logic;
signal bh3_w1_4 :  std_logic;
signal bh3_w2_4 :  std_logic;
signal bh3_w3_4 :  std_logic;
signal bh3_w4_4 :  std_logic;
signal bh3_w5_4 :  std_logic;
signal bh3_w6_4 :  std_logic;
signal bh3_w7_4 :  std_logic;
signal bh3_w8_4 :  std_logic;
signal bh3_w9_4 :  std_logic;
signal bh3_w10_4 :  std_logic;
signal bh3_w11_4 :  std_logic;
signal bh3_w12_4 :  std_logic;
signal bh3_w13_4 :  std_logic;
signal bh3_w14_4 :  std_logic;
signal bh3_w15_4 :  std_logic;
signal bh3_w16_4 :  std_logic;
signal bh3_w17_4 :  std_logic;
signal bh3_w18_4 :  std_logic;
signal bh3_w19_4 :  std_logic;
signal iX5 :  unsigned(19-0 downto 0);
signal bh3_w0_5 :  std_logic;
signal bh3_w1_5 :  std_logic;
signal bh3_w2_5 :  std_logic;
signal bh3_w3_5 :  std_logic;
signal bh3_w4_5 :  std_logic;
signal bh3_w5_5 :  std_logic;
signal bh3_w6_5 :  std_logic;
signal bh3_w7_5 :  std_logic;
signal bh3_w8_5 :  std_logic;
signal bh3_w9_5 :  std_logic;
signal bh3_w10_5 :  std_logic;
signal bh3_w11_5 :  std_logic;
signal bh3_w12_5 :  std_logic;
signal bh3_w13_5 :  std_logic;
signal bh3_w14_5 :  std_logic;
signal bh3_w15_5 :  std_logic;
signal bh3_w16_5 :  std_logic;
signal bh3_w17_5 :  std_logic;
signal bh3_w18_5 :  std_logic;
signal bh3_w19_5 :  std_logic;
signal iX6 :  unsigned(19-0 downto 0);
signal bh3_w0_6 :  std_logic;
signal bh3_w1_6 :  std_logic;
signal bh3_w2_6 :  std_logic;
signal bh3_w3_6 :  std_logic;
signal bh3_w4_6 :  std_logic;
signal bh3_w5_6 :  std_logic;
signal bh3_w6_6 :  std_logic;
signal bh3_w7_6 :  std_logic;
signal bh3_w8_6 :  std_logic;
signal bh3_w9_6 :  std_logic;
signal bh3_w10_6 :  std_logic;
signal bh3_w11_6 :  std_logic;
signal bh3_w12_6 :  std_logic;
signal bh3_w13_6 :  std_logic;
signal bh3_w14_6 :  std_logic;
signal bh3_w15_6 :  std_logic;
signal bh3_w16_6 :  std_logic;
signal bh3_w17_6 :  std_logic;
signal bh3_w18_6 :  std_logic;
signal bh3_w19_6 :  std_logic;
signal iX7 :  unsigned(19-0 downto 0);
signal bh3_w0_7 :  std_logic;
signal bh3_w1_7 :  std_logic;
signal bh3_w2_7 :  std_logic;
signal bh3_w3_7 :  std_logic;
signal bh3_w4_7 :  std_logic;
signal bh3_w5_7 :  std_logic;
signal bh3_w6_7 :  std_logic;
signal bh3_w7_7 :  std_logic;
signal bh3_w8_7 :  std_logic;
signal bh3_w9_7 :  std_logic;
signal bh3_w10_7 :  std_logic;
signal bh3_w11_7 :  std_logic;
signal bh3_w12_7 :  std_logic;
signal bh3_w13_7 :  std_logic;
signal bh3_w14_7 :  std_logic;
signal bh3_w15_7 :  std_logic;
signal bh3_w16_7 :  std_logic;
signal bh3_w17_7 :  std_logic;
signal bh3_w18_7 :  std_logic;
signal bh3_w19_7 :  std_logic;
signal iX8 :  unsigned(19-0 downto 0);
signal bh3_w0_8 :  std_logic;
signal bh3_w1_8 :  std_logic;
signal bh3_w2_8 :  std_logic;
signal bh3_w3_8 :  std_logic;
signal bh3_w4_8 :  std_logic;
signal bh3_w5_8 :  std_logic;
signal bh3_w6_8 :  std_logic;
signal bh3_w7_8 :  std_logic;
signal bh3_w8_8 :  std_logic;
signal bh3_w9_8 :  std_logic;
signal bh3_w10_8 :  std_logic;
signal bh3_w11_8 :  std_logic;
signal bh3_w12_8 :  std_logic;
signal bh3_w13_8 :  std_logic;
signal bh3_w14_8 :  std_logic;
signal bh3_w15_8 :  std_logic;
signal bh3_w16_8 :  std_logic;
signal bh3_w17_8 :  std_logic;
signal bh3_w18_8 :  std_logic;
signal bh3_w19_8 :  std_logic;
signal iX9 :  unsigned(19-0 downto 0);
signal bh3_w0_9 :  std_logic;
signal bh3_w1_9 :  std_logic;
signal bh3_w2_9 :  std_logic;
signal bh3_w3_9 :  std_logic;
signal bh3_w4_9 :  std_logic;
signal bh3_w5_9 :  std_logic;
signal bh3_w6_9 :  std_logic;
signal bh3_w7_9 :  std_logic;
signal bh3_w8_9 :  std_logic;
signal bh3_w9_9 :  std_logic;
signal bh3_w10_9 :  std_logic;
signal bh3_w11_9 :  std_logic;
signal bh3_w12_9 :  std_logic;
signal bh3_w13_9 :  std_logic;
signal bh3_w14_9 :  std_logic;
signal bh3_w15_9 :  std_logic;
signal bh3_w16_9 :  std_logic;
signal bh3_w17_9 :  std_logic;
signal bh3_w18_9 :  std_logic;
signal bh3_w19_9 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid7_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid7_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid7_Out0_copy8 :  std_logic_vector(2 downto 0);
signal bh3_w0_10 :  std_logic;
signal bh3_w1_10 :  std_logic;
signal bh3_w2_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid11_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid11_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid11_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid11_Out0_copy12 :  std_logic_vector(2 downto 0);
signal bh3_w0_11 :  std_logic;
signal bh3_w1_11 :  std_logic;
signal bh3_w2_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid13_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid13_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid13_Out0_copy14 :  std_logic_vector(2 downto 0);
signal bh3_w1_12 :  std_logic;
signal bh3_w2_12 :  std_logic;
signal bh3_w3_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid17_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid17_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid17_Out0_copy18 :  std_logic_vector(1 downto 0);
signal bh3_w1_13 :  std_logic;
signal bh3_w2_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid19_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid19_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid19_Out0_copy20 :  std_logic_vector(2 downto 0);
signal bh3_w2_14 :  std_logic;
signal bh3_w3_11 :  std_logic;
signal bh3_w4_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid21_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid21_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid21_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid21_Out0_copy22 :  std_logic_vector(2 downto 0);
signal bh3_w2_15 :  std_logic;
signal bh3_w3_12 :  std_logic;
signal bh3_w4_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid23_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid23_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid23_Out0_copy24 :  std_logic_vector(2 downto 0);
signal bh3_w3_13 :  std_logic;
signal bh3_w4_12 :  std_logic;
signal bh3_w5_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid25_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid25_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid25_Out0_copy26 :  std_logic_vector(1 downto 0);
signal bh3_w3_14 :  std_logic;
signal bh3_w4_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid27_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid27_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid27_Out0_copy28 :  std_logic_vector(2 downto 0);
signal bh3_w4_14 :  std_logic;
signal bh3_w5_11 :  std_logic;
signal bh3_w6_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid29_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid29_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid29_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid29_Out0_copy30 :  std_logic_vector(2 downto 0);
signal bh3_w4_15 :  std_logic;
signal bh3_w5_12 :  std_logic;
signal bh3_w6_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid31_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid31_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid31_Out0_copy32 :  std_logic_vector(2 downto 0);
signal bh3_w5_13 :  std_logic;
signal bh3_w6_12 :  std_logic;
signal bh3_w7_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid33_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid33_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid33_Out0_copy34 :  std_logic_vector(1 downto 0);
signal bh3_w5_14 :  std_logic;
signal bh3_w6_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid35_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid35_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid35_Out0_copy36 :  std_logic_vector(2 downto 0);
signal bh3_w6_14 :  std_logic;
signal bh3_w7_11 :  std_logic;
signal bh3_w8_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid37_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid37_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid37_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid37_Out0_copy38 :  std_logic_vector(2 downto 0);
signal bh3_w6_15 :  std_logic;
signal bh3_w7_12 :  std_logic;
signal bh3_w8_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid39_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid39_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid39_Out0_copy40 :  std_logic_vector(2 downto 0);
signal bh3_w7_13 :  std_logic;
signal bh3_w8_12 :  std_logic;
signal bh3_w9_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid41_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid41_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid41_Out0_copy42 :  std_logic_vector(1 downto 0);
signal bh3_w7_14 :  std_logic;
signal bh3_w8_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid43_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid43_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid43_Out0_copy44 :  std_logic_vector(2 downto 0);
signal bh3_w8_14 :  std_logic;
signal bh3_w9_11 :  std_logic;
signal bh3_w10_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid45_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid45_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid45_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid45_Out0_copy46 :  std_logic_vector(2 downto 0);
signal bh3_w8_15 :  std_logic;
signal bh3_w9_12 :  std_logic;
signal bh3_w10_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid47_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid47_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid47_Out0_copy48 :  std_logic_vector(2 downto 0);
signal bh3_w9_13 :  std_logic;
signal bh3_w10_12 :  std_logic;
signal bh3_w11_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid49_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid49_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid49_Out0_copy50 :  std_logic_vector(1 downto 0);
signal bh3_w9_14 :  std_logic;
signal bh3_w10_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid51_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid51_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid51_Out0_copy52 :  std_logic_vector(2 downto 0);
signal bh3_w10_14 :  std_logic;
signal bh3_w11_11 :  std_logic;
signal bh3_w12_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid53_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid53_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid53_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid53_Out0_copy54 :  std_logic_vector(2 downto 0);
signal bh3_w10_15 :  std_logic;
signal bh3_w11_12 :  std_logic;
signal bh3_w12_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid55_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid55_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid55_Out0_copy56 :  std_logic_vector(2 downto 0);
signal bh3_w11_13 :  std_logic;
signal bh3_w12_12 :  std_logic;
signal bh3_w13_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid57_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid57_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid57_Out0_copy58 :  std_logic_vector(1 downto 0);
signal bh3_w11_14 :  std_logic;
signal bh3_w12_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid59_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid59_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid59_Out0_copy60 :  std_logic_vector(2 downto 0);
signal bh3_w12_14 :  std_logic;
signal bh3_w13_11 :  std_logic;
signal bh3_w14_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid61_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid61_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid61_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid61_Out0_copy62 :  std_logic_vector(2 downto 0);
signal bh3_w12_15 :  std_logic;
signal bh3_w13_12 :  std_logic;
signal bh3_w14_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid63_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid63_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid63_Out0_copy64 :  std_logic_vector(2 downto 0);
signal bh3_w13_13 :  std_logic;
signal bh3_w14_12 :  std_logic;
signal bh3_w15_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid65_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid65_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid65_Out0_copy66 :  std_logic_vector(1 downto 0);
signal bh3_w13_14 :  std_logic;
signal bh3_w14_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid67_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid67_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid67_Out0_copy68 :  std_logic_vector(2 downto 0);
signal bh3_w14_14 :  std_logic;
signal bh3_w15_11 :  std_logic;
signal bh3_w16_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid69_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid69_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid69_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid69_Out0_copy70 :  std_logic_vector(2 downto 0);
signal bh3_w14_15 :  std_logic;
signal bh3_w15_12 :  std_logic;
signal bh3_w16_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid71_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid71_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid71_Out0_copy72 :  std_logic_vector(2 downto 0);
signal bh3_w15_13 :  std_logic;
signal bh3_w16_12 :  std_logic;
signal bh3_w17_10 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid73_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid73_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid73_Out0_copy74 :  std_logic_vector(1 downto 0);
signal bh3_w15_14 :  std_logic;
signal bh3_w16_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid75_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid75_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid75_Out0_copy76 :  std_logic_vector(2 downto 0);
signal bh3_w16_14 :  std_logic;
signal bh3_w17_11 :  std_logic;
signal bh3_w18_10 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid77_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid77_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid77_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid77_Out0_copy78 :  std_logic_vector(2 downto 0);
signal bh3_w16_15 :  std_logic;
signal bh3_w17_12 :  std_logic;
signal bh3_w18_11 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid79_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid79_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid79_Out0_copy80 :  std_logic_vector(2 downto 0);
signal bh3_w17_13 :  std_logic;
signal bh3_w18_12 :  std_logic;
signal bh3_w19_10, bh3_w19_10_d1 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid81_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid81_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid81_Out0_copy82 :  std_logic_vector(1 downto 0);
signal bh3_w17_14 :  std_logic;
signal bh3_w18_13 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid83_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid83_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid83_Out0_copy84 :  std_logic_vector(2 downto 0);
signal bh3_w18_14 :  std_logic;
signal bh3_w19_11 :  std_logic;
signal bh3_w20_0 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid85_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid85_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid85_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid85_Out0_copy86 :  std_logic_vector(2 downto 0);
signal bh3_w18_15 :  std_logic;
signal bh3_w19_12 :  std_logic;
signal bh3_w20_1 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid87_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid87_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid87_Out0_copy88 :  std_logic_vector(2 downto 0);
signal bh3_w19_13 :  std_logic;
signal bh3_w20_2 :  std_logic;
signal bh3_w21_0, bh3_w21_0_d1 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid89_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid89_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid89_Out0_copy90 :  std_logic_vector(1 downto 0);
signal bh3_w19_14 :  std_logic;
signal bh3_w20_3 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid91_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid91_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid91_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92, Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92_d1 :  std_logic_vector(2 downto 0);
signal bh3_w0_12 :  std_logic;
signal bh3_w1_14 :  std_logic;
signal bh3_w2_16 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid93_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid93_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94, Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94_d1 :  std_logic_vector(1 downto 0);
signal bh3_w1_15 :  std_logic;
signal bh3_w2_17 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid95_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid95_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96, Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96_d1 :  std_logic_vector(2 downto 0);
signal bh3_w2_18 :  std_logic;
signal bh3_w3_15 :  std_logic;
signal bh3_w4_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid99_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid99_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100, Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100_d1 :  std_logic_vector(2 downto 0);
signal bh3_w3_16 :  std_logic;
signal bh3_w4_17 :  std_logic;
signal bh3_w5_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid101_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid101_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102, Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102_d1 :  std_logic_vector(2 downto 0);
signal bh3_w4_18 :  std_logic;
signal bh3_w5_16 :  std_logic;
signal bh3_w6_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid103_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid103_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104, Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104_d1 :  std_logic_vector(2 downto 0);
signal bh3_w5_17 :  std_logic;
signal bh3_w6_17 :  std_logic;
signal bh3_w7_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid105_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid105_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106, Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106_d1 :  std_logic_vector(2 downto 0);
signal bh3_w6_18 :  std_logic;
signal bh3_w7_16 :  std_logic;
signal bh3_w8_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid107_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid107_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108, Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108_d1 :  std_logic_vector(2 downto 0);
signal bh3_w7_17 :  std_logic;
signal bh3_w8_17 :  std_logic;
signal bh3_w9_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid109_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid109_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110, Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110_d1 :  std_logic_vector(2 downto 0);
signal bh3_w8_18 :  std_logic;
signal bh3_w9_16 :  std_logic;
signal bh3_w10_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid111_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid111_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112, Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112_d1 :  std_logic_vector(2 downto 0);
signal bh3_w9_17 :  std_logic;
signal bh3_w10_17 :  std_logic;
signal bh3_w11_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid113_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid113_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114, Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114_d1 :  std_logic_vector(2 downto 0);
signal bh3_w10_18 :  std_logic;
signal bh3_w11_16 :  std_logic;
signal bh3_w12_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid115_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid115_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116, Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116_d1 :  std_logic_vector(2 downto 0);
signal bh3_w11_17 :  std_logic;
signal bh3_w12_17 :  std_logic;
signal bh3_w13_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid117_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid117_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118, Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118_d1 :  std_logic_vector(2 downto 0);
signal bh3_w12_18 :  std_logic;
signal bh3_w13_16 :  std_logic;
signal bh3_w14_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid119_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid119_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120, Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120_d1 :  std_logic_vector(2 downto 0);
signal bh3_w13_17 :  std_logic;
signal bh3_w14_17 :  std_logic;
signal bh3_w15_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid121_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid121_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122, Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122_d1 :  std_logic_vector(2 downto 0);
signal bh3_w14_18 :  std_logic;
signal bh3_w15_16 :  std_logic;
signal bh3_w16_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid123_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid123_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124, Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124_d1 :  std_logic_vector(2 downto 0);
signal bh3_w15_17 :  std_logic;
signal bh3_w16_17 :  std_logic;
signal bh3_w17_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid125_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid125_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126, Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126_d1 :  std_logic_vector(2 downto 0);
signal bh3_w16_18 :  std_logic;
signal bh3_w17_16 :  std_logic;
signal bh3_w18_16 :  std_logic;
signal Compressor_5_3_F800_uid98_bh3_uid127_In0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid127_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128, Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128_d1 :  std_logic_vector(2 downto 0);
signal bh3_w17_17 :  std_logic;
signal bh3_w18_17 :  std_logic;
signal bh3_w19_15 :  std_logic;
signal Compressor_6_3_F800_uid6_bh3_uid129_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid129_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130, Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130_d1 :  std_logic_vector(2 downto 0);
signal bh3_w18_18 :  std_logic;
signal bh3_w19_16 :  std_logic;
signal bh3_w20_4 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid131_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid131_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid131_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132, Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132_d1 :  std_logic_vector(2 downto 0);
signal bh3_w19_17 :  std_logic;
signal bh3_w20_5 :  std_logic;
signal bh3_w21_1 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid133_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid133_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134, Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134_d1 :  std_logic_vector(1 downto 0);
signal bh3_w20_6 :  std_logic;
signal bh3_w21_2 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid137_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid137_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid137_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid137_Out0_copy138 :  std_logic_vector(2 downto 0);
signal bh3_w0_13, bh3_w0_13_d1 :  std_logic;
signal bh3_w1_16, bh3_w1_16_d1 :  std_logic;
signal bh3_w2_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid139_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid139_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid139_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid139_Out0_copy140 :  std_logic_vector(2 downto 0);
signal bh3_w2_20 :  std_logic;
signal bh3_w3_17 :  std_logic;
signal bh3_w4_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid141_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid141_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid141_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid141_Out0_copy142 :  std_logic_vector(2 downto 0);
signal bh3_w4_20 :  std_logic;
signal bh3_w5_18 :  std_logic;
signal bh3_w6_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid143_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid143_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid143_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid143_Out0_copy144 :  std_logic_vector(2 downto 0);
signal bh3_w6_20 :  std_logic;
signal bh3_w7_18 :  std_logic;
signal bh3_w8_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid145_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid145_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid145_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid145_Out0_copy146 :  std_logic_vector(2 downto 0);
signal bh3_w8_20 :  std_logic;
signal bh3_w9_18 :  std_logic;
signal bh3_w10_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid147_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid147_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid147_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid147_Out0_copy148 :  std_logic_vector(2 downto 0);
signal bh3_w10_20 :  std_logic;
signal bh3_w11_18 :  std_logic;
signal bh3_w12_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid149_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid149_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid149_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid149_Out0_copy150 :  std_logic_vector(2 downto 0);
signal bh3_w12_20 :  std_logic;
signal bh3_w13_18 :  std_logic;
signal bh3_w14_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid151_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid151_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid151_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid151_Out0_copy152 :  std_logic_vector(2 downto 0);
signal bh3_w14_20 :  std_logic;
signal bh3_w15_18 :  std_logic;
signal bh3_w16_19 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid153_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid153_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid153_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid153_Out0_copy154 :  std_logic_vector(2 downto 0);
signal bh3_w16_20 :  std_logic;
signal bh3_w17_18 :  std_logic;
signal bh3_w18_19 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid155_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid155_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid155_Out0_copy156 :  std_logic_vector(1 downto 0);
signal bh3_w18_20 :  std_logic;
signal bh3_w19_18 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid157_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid157_In1, Compressor_14_3_F800_uid10_bh3_uid157_In1_d1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid157_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid157_Out0_copy158 :  std_logic_vector(2 downto 0);
signal bh3_w19_19 :  std_logic;
signal bh3_w20_7 :  std_logic;
signal bh3_w21_3 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid159_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid159_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid159_Out0_copy160 :  std_logic_vector(1 downto 0);
signal bh3_w20_8 :  std_logic;
signal bh3_w21_4 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid161_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid161_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid161_Out0_copy162 :  std_logic_vector(1 downto 0);
signal bh3_w21_5 :  std_logic;
signal bh3_w22_0, bh3_w22_0_d1 :  std_logic;
signal Compressor_14_3_F800_uid10_bh3_uid163_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid163_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid163_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164, Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164_d1 :  std_logic_vector(2 downto 0);
signal bh3_w2_21 :  std_logic;
signal bh3_w3_18 :  std_logic;
signal bh3_w4_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid165_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid165_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid165_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166, Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166_d1 :  std_logic_vector(2 downto 0);
signal bh3_w4_22 :  std_logic;
signal bh3_w5_19 :  std_logic;
signal bh3_w6_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid167_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid167_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid167_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168, Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168_d1 :  std_logic_vector(2 downto 0);
signal bh3_w6_22 :  std_logic;
signal bh3_w7_19 :  std_logic;
signal bh3_w8_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid169_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid169_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid169_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170, Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170_d1 :  std_logic_vector(2 downto 0);
signal bh3_w8_22 :  std_logic;
signal bh3_w9_19 :  std_logic;
signal bh3_w10_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid171_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid171_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid171_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172, Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172_d1 :  std_logic_vector(2 downto 0);
signal bh3_w10_22 :  std_logic;
signal bh3_w11_19 :  std_logic;
signal bh3_w12_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid173_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid173_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid173_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174, Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174_d1 :  std_logic_vector(2 downto 0);
signal bh3_w12_22 :  std_logic;
signal bh3_w13_19 :  std_logic;
signal bh3_w14_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid175_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid175_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid175_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176, Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176_d1 :  std_logic_vector(2 downto 0);
signal bh3_w14_22 :  std_logic;
signal bh3_w15_19 :  std_logic;
signal bh3_w16_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid177_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid177_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid177_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178, Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178_d1 :  std_logic_vector(2 downto 0);
signal bh3_w16_22 :  std_logic;
signal bh3_w17_19 :  std_logic;
signal bh3_w18_21 :  std_logic;
signal Compressor_23_3_F800_uid136_bh3_uid179_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid179_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid179_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180, Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180_d1 :  std_logic_vector(2 downto 0);
signal bh3_w18_22 :  std_logic;
signal bh3_w19_20 :  std_logic;
signal bh3_w20_9 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid181_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid181_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182, Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182_d1 :  std_logic_vector(1 downto 0);
signal bh3_w20_10 :  std_logic;
signal bh3_w21_6 :  std_logic;
signal Compressor_3_2_F800_uid16_bh3_uid183_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid183_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184, Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184_d1 :  std_logic_vector(1 downto 0);
signal bh3_w21_7 :  std_logic;
signal bh3_w22_1 :  std_logic;
signal tmp_bitheapResult_bh3_3, tmp_bitheapResult_bh3_3_d1, tmp_bitheapResult_bh3_3_d2 :  std_logic_vector(3 downto 0);
signal bitheapFinalAdd_bh3_In0 :  std_logic_vector(20 downto 0);
signal bitheapFinalAdd_bh3_In1 :  std_logic_vector(20 downto 0);
signal bitheapFinalAdd_bh3_Cin :  std_logic;
signal bitheapFinalAdd_bh3_Out :  std_logic_vector(20 downto 0);
signal bitheapResult_bh3 :  std_logic_vector(23 downto 0);
signal OutRes :  std_logic_vector(23 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            bh3_w19_10_d1 <=  bh3_w19_10;
            bh3_w21_0_d1 <=  bh3_w21_0;
            Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92_d1 <=  Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92;
            Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94_d1 <=  Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94;
            Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96_d1 <=  Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96;
            Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100_d1 <=  Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100;
            Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102_d1 <=  Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102;
            Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104_d1 <=  Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104;
            Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106_d1 <=  Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106;
            Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108_d1 <=  Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108;
            Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110_d1 <=  Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110;
            Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112_d1 <=  Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112;
            Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114_d1 <=  Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114;
            Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116_d1 <=  Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116;
            Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118_d1 <=  Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118;
            Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120_d1 <=  Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120;
            Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122_d1 <=  Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122;
            Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124_d1 <=  Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124;
            Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126_d1 <=  Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126;
            Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128_d1 <=  Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128;
            Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130_d1 <=  Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130;
            Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132_d1 <=  Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132;
            Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134_d1 <=  Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134;
            bh3_w0_13_d1 <=  bh3_w0_13;
            bh3_w1_16_d1 <=  bh3_w1_16;
            Compressor_14_3_F800_uid10_bh3_uid157_In1_d1 <=  Compressor_14_3_F800_uid10_bh3_uid157_In1;
            bh3_w22_0_d1 <=  bh3_w22_0;
            Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164_d1 <=  Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164;
            Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166_d1 <=  Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166;
            Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168_d1 <=  Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168;
            Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170_d1 <=  Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170;
            Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172_d1 <=  Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172;
            Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174_d1 <=  Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174;
            Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176_d1 <=  Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176;
            Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178_d1 <=  Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178;
            Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180_d1 <=  Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180;
            Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182_d1 <=  Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182;
            Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184_d1 <=  Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184;
            tmp_bitheapResult_bh3_3_d1 <=  tmp_bitheapResult_bh3_3;
            tmp_bitheapResult_bh3_3_d2 <=  tmp_bitheapResult_bh3_3_d1;
         end if;
      end process;
   iX0 <= unsigned(X0);
   bh3_w0_0 <= iX0(0);
   bh3_w1_0 <= iX0(1);
   bh3_w2_0 <= iX0(2);
   bh3_w3_0 <= iX0(3);
   bh3_w4_0 <= iX0(4);
   bh3_w5_0 <= iX0(5);
   bh3_w6_0 <= iX0(6);
   bh3_w7_0 <= iX0(7);
   bh3_w8_0 <= iX0(8);
   bh3_w9_0 <= iX0(9);
   bh3_w10_0 <= iX0(10);
   bh3_w11_0 <= iX0(11);
   bh3_w12_0 <= iX0(12);
   bh3_w13_0 <= iX0(13);
   bh3_w14_0 <= iX0(14);
   bh3_w15_0 <= iX0(15);
   bh3_w16_0 <= iX0(16);
   bh3_w17_0 <= iX0(17);
   bh3_w18_0 <= iX0(18);
   bh3_w19_0 <= iX0(19);
   iX1 <= unsigned(X1);
   bh3_w0_1 <= iX1(0);
   bh3_w1_1 <= iX1(1);
   bh3_w2_1 <= iX1(2);
   bh3_w3_1 <= iX1(3);
   bh3_w4_1 <= iX1(4);
   bh3_w5_1 <= iX1(5);
   bh3_w6_1 <= iX1(6);
   bh3_w7_1 <= iX1(7);
   bh3_w8_1 <= iX1(8);
   bh3_w9_1 <= iX1(9);
   bh3_w10_1 <= iX1(10);
   bh3_w11_1 <= iX1(11);
   bh3_w12_1 <= iX1(12);
   bh3_w13_1 <= iX1(13);
   bh3_w14_1 <= iX1(14);
   bh3_w15_1 <= iX1(15);
   bh3_w16_1 <= iX1(16);
   bh3_w17_1 <= iX1(17);
   bh3_w18_1 <= iX1(18);
   bh3_w19_1 <= iX1(19);
   iX2 <= unsigned(X2);
   bh3_w0_2 <= iX2(0);
   bh3_w1_2 <= iX2(1);
   bh3_w2_2 <= iX2(2);
   bh3_w3_2 <= iX2(3);
   bh3_w4_2 <= iX2(4);
   bh3_w5_2 <= iX2(5);
   bh3_w6_2 <= iX2(6);
   bh3_w7_2 <= iX2(7);
   bh3_w8_2 <= iX2(8);
   bh3_w9_2 <= iX2(9);
   bh3_w10_2 <= iX2(10);
   bh3_w11_2 <= iX2(11);
   bh3_w12_2 <= iX2(12);
   bh3_w13_2 <= iX2(13);
   bh3_w14_2 <= iX2(14);
   bh3_w15_2 <= iX2(15);
   bh3_w16_2 <= iX2(16);
   bh3_w17_2 <= iX2(17);
   bh3_w18_2 <= iX2(18);
   bh3_w19_2 <= iX2(19);
   iX3 <= unsigned(X3);
   bh3_w0_3 <= iX3(0);
   bh3_w1_3 <= iX3(1);
   bh3_w2_3 <= iX3(2);
   bh3_w3_3 <= iX3(3);
   bh3_w4_3 <= iX3(4);
   bh3_w5_3 <= iX3(5);
   bh3_w6_3 <= iX3(6);
   bh3_w7_3 <= iX3(7);
   bh3_w8_3 <= iX3(8);
   bh3_w9_3 <= iX3(9);
   bh3_w10_3 <= iX3(10);
   bh3_w11_3 <= iX3(11);
   bh3_w12_3 <= iX3(12);
   bh3_w13_3 <= iX3(13);
   bh3_w14_3 <= iX3(14);
   bh3_w15_3 <= iX3(15);
   bh3_w16_3 <= iX3(16);
   bh3_w17_3 <= iX3(17);
   bh3_w18_3 <= iX3(18);
   bh3_w19_3 <= iX3(19);
   iX4 <= unsigned(X4);
   bh3_w0_4 <= iX4(0);
   bh3_w1_4 <= iX4(1);
   bh3_w2_4 <= iX4(2);
   bh3_w3_4 <= iX4(3);
   bh3_w4_4 <= iX4(4);
   bh3_w5_4 <= iX4(5);
   bh3_w6_4 <= iX4(6);
   bh3_w7_4 <= iX4(7);
   bh3_w8_4 <= iX4(8);
   bh3_w9_4 <= iX4(9);
   bh3_w10_4 <= iX4(10);
   bh3_w11_4 <= iX4(11);
   bh3_w12_4 <= iX4(12);
   bh3_w13_4 <= iX4(13);
   bh3_w14_4 <= iX4(14);
   bh3_w15_4 <= iX4(15);
   bh3_w16_4 <= iX4(16);
   bh3_w17_4 <= iX4(17);
   bh3_w18_4 <= iX4(18);
   bh3_w19_4 <= iX4(19);
   iX5 <= unsigned(X5);
   bh3_w0_5 <= iX5(0);
   bh3_w1_5 <= iX5(1);
   bh3_w2_5 <= iX5(2);
   bh3_w3_5 <= iX5(3);
   bh3_w4_5 <= iX5(4);
   bh3_w5_5 <= iX5(5);
   bh3_w6_5 <= iX5(6);
   bh3_w7_5 <= iX5(7);
   bh3_w8_5 <= iX5(8);
   bh3_w9_5 <= iX5(9);
   bh3_w10_5 <= iX5(10);
   bh3_w11_5 <= iX5(11);
   bh3_w12_5 <= iX5(12);
   bh3_w13_5 <= iX5(13);
   bh3_w14_5 <= iX5(14);
   bh3_w15_5 <= iX5(15);
   bh3_w16_5 <= iX5(16);
   bh3_w17_5 <= iX5(17);
   bh3_w18_5 <= iX5(18);
   bh3_w19_5 <= iX5(19);
   iX6 <= unsigned(X6);
   bh3_w0_6 <= iX6(0);
   bh3_w1_6 <= iX6(1);
   bh3_w2_6 <= iX6(2);
   bh3_w3_6 <= iX6(3);
   bh3_w4_6 <= iX6(4);
   bh3_w5_6 <= iX6(5);
   bh3_w6_6 <= iX6(6);
   bh3_w7_6 <= iX6(7);
   bh3_w8_6 <= iX6(8);
   bh3_w9_6 <= iX6(9);
   bh3_w10_6 <= iX6(10);
   bh3_w11_6 <= iX6(11);
   bh3_w12_6 <= iX6(12);
   bh3_w13_6 <= iX6(13);
   bh3_w14_6 <= iX6(14);
   bh3_w15_6 <= iX6(15);
   bh3_w16_6 <= iX6(16);
   bh3_w17_6 <= iX6(17);
   bh3_w18_6 <= iX6(18);
   bh3_w19_6 <= iX6(19);
   iX7 <= unsigned(X7);
   bh3_w0_7 <= iX7(0);
   bh3_w1_7 <= iX7(1);
   bh3_w2_7 <= iX7(2);
   bh3_w3_7 <= iX7(3);
   bh3_w4_7 <= iX7(4);
   bh3_w5_7 <= iX7(5);
   bh3_w6_7 <= iX7(6);
   bh3_w7_7 <= iX7(7);
   bh3_w8_7 <= iX7(8);
   bh3_w9_7 <= iX7(9);
   bh3_w10_7 <= iX7(10);
   bh3_w11_7 <= iX7(11);
   bh3_w12_7 <= iX7(12);
   bh3_w13_7 <= iX7(13);
   bh3_w14_7 <= iX7(14);
   bh3_w15_7 <= iX7(15);
   bh3_w16_7 <= iX7(16);
   bh3_w17_7 <= iX7(17);
   bh3_w18_7 <= iX7(18);
   bh3_w19_7 <= iX7(19);
   iX8 <= unsigned(X8);
   bh3_w0_8 <= iX8(0);
   bh3_w1_8 <= iX8(1);
   bh3_w2_8 <= iX8(2);
   bh3_w3_8 <= iX8(3);
   bh3_w4_8 <= iX8(4);
   bh3_w5_8 <= iX8(5);
   bh3_w6_8 <= iX8(6);
   bh3_w7_8 <= iX8(7);
   bh3_w8_8 <= iX8(8);
   bh3_w9_8 <= iX8(9);
   bh3_w10_8 <= iX8(10);
   bh3_w11_8 <= iX8(11);
   bh3_w12_8 <= iX8(12);
   bh3_w13_8 <= iX8(13);
   bh3_w14_8 <= iX8(14);
   bh3_w15_8 <= iX8(15);
   bh3_w16_8 <= iX8(16);
   bh3_w17_8 <= iX8(17);
   bh3_w18_8 <= iX8(18);
   bh3_w19_8 <= iX8(19);
   iX9 <= unsigned(X9);
   bh3_w0_9 <= iX9(0);
   bh3_w1_9 <= iX9(1);
   bh3_w2_9 <= iX9(2);
   bh3_w3_9 <= iX9(3);
   bh3_w4_9 <= iX9(4);
   bh3_w5_9 <= iX9(5);
   bh3_w6_9 <= iX9(6);
   bh3_w7_9 <= iX9(7);
   bh3_w8_9 <= iX9(8);
   bh3_w9_9 <= iX9(9);
   bh3_w10_9 <= iX9(10);
   bh3_w11_9 <= iX9(11);
   bh3_w12_9 <= iX9(12);
   bh3_w13_9 <= iX9(13);
   bh3_w14_9 <= iX9(14);
   bh3_w15_9 <= iX9(15);
   bh3_w16_9 <= iX9(16);
   bh3_w17_9 <= iX9(17);
   bh3_w18_9 <= iX9(18);
   bh3_w19_9 <= iX9(19);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_6_3_F800_uid6_bh3_uid7_In0 <= "" & bh3_w0_0 & bh3_w0_1 & bh3_w0_2 & bh3_w0_3 & bh3_w0_4 & bh3_w0_5;
   Compressor_6_3_F800_uid6_uid7: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid7_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid7_Out0_copy8);
   Compressor_6_3_F800_uid6_bh3_uid7_Out0 <= Compressor_6_3_F800_uid6_bh3_uid7_Out0_copy8; -- output copy to hold a pipeline register if needed

   bh3_w0_10 <= Compressor_6_3_F800_uid6_bh3_uid7_Out0(0);
   bh3_w1_10 <= Compressor_6_3_F800_uid6_bh3_uid7_Out0(1);
   bh3_w2_10 <= Compressor_6_3_F800_uid6_bh3_uid7_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid11_In0 <= "" & bh3_w0_6 & bh3_w0_7 & bh3_w0_8 & bh3_w0_9;
   Compressor_14_3_F800_uid10_bh3_uid11_In1 <= "" & bh3_w1_0;
   Compressor_14_3_F800_uid10_uid11: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid11_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid11_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid11_Out0_copy12);
   Compressor_14_3_F800_uid10_bh3_uid11_Out0 <= Compressor_14_3_F800_uid10_bh3_uid11_Out0_copy12; -- output copy to hold a pipeline register if needed

   bh3_w0_11 <= Compressor_14_3_F800_uid10_bh3_uid11_Out0(0);
   bh3_w1_11 <= Compressor_14_3_F800_uid10_bh3_uid11_Out0(1);
   bh3_w2_11 <= Compressor_14_3_F800_uid10_bh3_uid11_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid13_In0 <= "" & bh3_w1_1 & bh3_w1_2 & bh3_w1_3 & bh3_w1_4 & bh3_w1_5 & bh3_w1_6;
   Compressor_6_3_F800_uid6_uid13: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid13_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid13_Out0_copy14);
   Compressor_6_3_F800_uid6_bh3_uid13_Out0 <= Compressor_6_3_F800_uid6_bh3_uid13_Out0_copy14; -- output copy to hold a pipeline register if needed

   bh3_w1_12 <= Compressor_6_3_F800_uid6_bh3_uid13_Out0(0);
   bh3_w2_12 <= Compressor_6_3_F800_uid6_bh3_uid13_Out0(1);
   bh3_w3_10 <= Compressor_6_3_F800_uid6_bh3_uid13_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid17_In0 <= "" & bh3_w1_7 & bh3_w1_8 & bh3_w1_9;
   Compressor_3_2_F800_uid16_uid17: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid17_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid17_Out0_copy18);
   Compressor_3_2_F800_uid16_bh3_uid17_Out0 <= Compressor_3_2_F800_uid16_bh3_uid17_Out0_copy18; -- output copy to hold a pipeline register if needed

   bh3_w1_13 <= Compressor_3_2_F800_uid16_bh3_uid17_Out0(0);
   bh3_w2_13 <= Compressor_3_2_F800_uid16_bh3_uid17_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid19_In0 <= "" & bh3_w2_0 & bh3_w2_1 & bh3_w2_2 & bh3_w2_3 & bh3_w2_4 & bh3_w2_5;
   Compressor_6_3_F800_uid6_uid19: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid19_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid19_Out0_copy20);
   Compressor_6_3_F800_uid6_bh3_uid19_Out0 <= Compressor_6_3_F800_uid6_bh3_uid19_Out0_copy20; -- output copy to hold a pipeline register if needed

   bh3_w2_14 <= Compressor_6_3_F800_uid6_bh3_uid19_Out0(0);
   bh3_w3_11 <= Compressor_6_3_F800_uid6_bh3_uid19_Out0(1);
   bh3_w4_10 <= Compressor_6_3_F800_uid6_bh3_uid19_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid21_In0 <= "" & bh3_w2_6 & bh3_w2_7 & bh3_w2_8 & bh3_w2_9;
   Compressor_14_3_F800_uid10_bh3_uid21_In1 <= "" & bh3_w3_0;
   Compressor_14_3_F800_uid10_uid21: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid21_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid21_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid21_Out0_copy22);
   Compressor_14_3_F800_uid10_bh3_uid21_Out0 <= Compressor_14_3_F800_uid10_bh3_uid21_Out0_copy22; -- output copy to hold a pipeline register if needed

   bh3_w2_15 <= Compressor_14_3_F800_uid10_bh3_uid21_Out0(0);
   bh3_w3_12 <= Compressor_14_3_F800_uid10_bh3_uid21_Out0(1);
   bh3_w4_11 <= Compressor_14_3_F800_uid10_bh3_uid21_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid23_In0 <= "" & bh3_w3_1 & bh3_w3_2 & bh3_w3_3 & bh3_w3_4 & bh3_w3_5 & bh3_w3_6;
   Compressor_6_3_F800_uid6_uid23: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid23_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid23_Out0_copy24);
   Compressor_6_3_F800_uid6_bh3_uid23_Out0 <= Compressor_6_3_F800_uid6_bh3_uid23_Out0_copy24; -- output copy to hold a pipeline register if needed

   bh3_w3_13 <= Compressor_6_3_F800_uid6_bh3_uid23_Out0(0);
   bh3_w4_12 <= Compressor_6_3_F800_uid6_bh3_uid23_Out0(1);
   bh3_w5_10 <= Compressor_6_3_F800_uid6_bh3_uid23_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid25_In0 <= "" & bh3_w3_7 & bh3_w3_8 & bh3_w3_9;
   Compressor_3_2_F800_uid16_uid25: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid25_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid25_Out0_copy26);
   Compressor_3_2_F800_uid16_bh3_uid25_Out0 <= Compressor_3_2_F800_uid16_bh3_uid25_Out0_copy26; -- output copy to hold a pipeline register if needed

   bh3_w3_14 <= Compressor_3_2_F800_uid16_bh3_uid25_Out0(0);
   bh3_w4_13 <= Compressor_3_2_F800_uid16_bh3_uid25_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid27_In0 <= "" & bh3_w4_0 & bh3_w4_1 & bh3_w4_2 & bh3_w4_3 & bh3_w4_4 & bh3_w4_5;
   Compressor_6_3_F800_uid6_uid27: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid27_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid27_Out0_copy28);
   Compressor_6_3_F800_uid6_bh3_uid27_Out0 <= Compressor_6_3_F800_uid6_bh3_uid27_Out0_copy28; -- output copy to hold a pipeline register if needed

   bh3_w4_14 <= Compressor_6_3_F800_uid6_bh3_uid27_Out0(0);
   bh3_w5_11 <= Compressor_6_3_F800_uid6_bh3_uid27_Out0(1);
   bh3_w6_10 <= Compressor_6_3_F800_uid6_bh3_uid27_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid29_In0 <= "" & bh3_w4_6 & bh3_w4_7 & bh3_w4_8 & bh3_w4_9;
   Compressor_14_3_F800_uid10_bh3_uid29_In1 <= "" & bh3_w5_0;
   Compressor_14_3_F800_uid10_uid29: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid29_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid29_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid29_Out0_copy30);
   Compressor_14_3_F800_uid10_bh3_uid29_Out0 <= Compressor_14_3_F800_uid10_bh3_uid29_Out0_copy30; -- output copy to hold a pipeline register if needed

   bh3_w4_15 <= Compressor_14_3_F800_uid10_bh3_uid29_Out0(0);
   bh3_w5_12 <= Compressor_14_3_F800_uid10_bh3_uid29_Out0(1);
   bh3_w6_11 <= Compressor_14_3_F800_uid10_bh3_uid29_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid31_In0 <= "" & bh3_w5_1 & bh3_w5_2 & bh3_w5_3 & bh3_w5_4 & bh3_w5_5 & bh3_w5_6;
   Compressor_6_3_F800_uid6_uid31: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid31_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid31_Out0_copy32);
   Compressor_6_3_F800_uid6_bh3_uid31_Out0 <= Compressor_6_3_F800_uid6_bh3_uid31_Out0_copy32; -- output copy to hold a pipeline register if needed

   bh3_w5_13 <= Compressor_6_3_F800_uid6_bh3_uid31_Out0(0);
   bh3_w6_12 <= Compressor_6_3_F800_uid6_bh3_uid31_Out0(1);
   bh3_w7_10 <= Compressor_6_3_F800_uid6_bh3_uid31_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid33_In0 <= "" & bh3_w5_7 & bh3_w5_8 & bh3_w5_9;
   Compressor_3_2_F800_uid16_uid33: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid33_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid33_Out0_copy34);
   Compressor_3_2_F800_uid16_bh3_uid33_Out0 <= Compressor_3_2_F800_uid16_bh3_uid33_Out0_copy34; -- output copy to hold a pipeline register if needed

   bh3_w5_14 <= Compressor_3_2_F800_uid16_bh3_uid33_Out0(0);
   bh3_w6_13 <= Compressor_3_2_F800_uid16_bh3_uid33_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid35_In0 <= "" & bh3_w6_0 & bh3_w6_1 & bh3_w6_2 & bh3_w6_3 & bh3_w6_4 & bh3_w6_5;
   Compressor_6_3_F800_uid6_uid35: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid35_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid35_Out0_copy36);
   Compressor_6_3_F800_uid6_bh3_uid35_Out0 <= Compressor_6_3_F800_uid6_bh3_uid35_Out0_copy36; -- output copy to hold a pipeline register if needed

   bh3_w6_14 <= Compressor_6_3_F800_uid6_bh3_uid35_Out0(0);
   bh3_w7_11 <= Compressor_6_3_F800_uid6_bh3_uid35_Out0(1);
   bh3_w8_10 <= Compressor_6_3_F800_uid6_bh3_uid35_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid37_In0 <= "" & bh3_w6_6 & bh3_w6_7 & bh3_w6_8 & bh3_w6_9;
   Compressor_14_3_F800_uid10_bh3_uid37_In1 <= "" & bh3_w7_0;
   Compressor_14_3_F800_uid10_uid37: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid37_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid37_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid37_Out0_copy38);
   Compressor_14_3_F800_uid10_bh3_uid37_Out0 <= Compressor_14_3_F800_uid10_bh3_uid37_Out0_copy38; -- output copy to hold a pipeline register if needed

   bh3_w6_15 <= Compressor_14_3_F800_uid10_bh3_uid37_Out0(0);
   bh3_w7_12 <= Compressor_14_3_F800_uid10_bh3_uid37_Out0(1);
   bh3_w8_11 <= Compressor_14_3_F800_uid10_bh3_uid37_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid39_In0 <= "" & bh3_w7_1 & bh3_w7_2 & bh3_w7_3 & bh3_w7_4 & bh3_w7_5 & bh3_w7_6;
   Compressor_6_3_F800_uid6_uid39: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid39_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid39_Out0_copy40);
   Compressor_6_3_F800_uid6_bh3_uid39_Out0 <= Compressor_6_3_F800_uid6_bh3_uid39_Out0_copy40; -- output copy to hold a pipeline register if needed

   bh3_w7_13 <= Compressor_6_3_F800_uid6_bh3_uid39_Out0(0);
   bh3_w8_12 <= Compressor_6_3_F800_uid6_bh3_uid39_Out0(1);
   bh3_w9_10 <= Compressor_6_3_F800_uid6_bh3_uid39_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid41_In0 <= "" & bh3_w7_7 & bh3_w7_8 & bh3_w7_9;
   Compressor_3_2_F800_uid16_uid41: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid41_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid41_Out0_copy42);
   Compressor_3_2_F800_uid16_bh3_uid41_Out0 <= Compressor_3_2_F800_uid16_bh3_uid41_Out0_copy42; -- output copy to hold a pipeline register if needed

   bh3_w7_14 <= Compressor_3_2_F800_uid16_bh3_uid41_Out0(0);
   bh3_w8_13 <= Compressor_3_2_F800_uid16_bh3_uid41_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid43_In0 <= "" & bh3_w8_0 & bh3_w8_1 & bh3_w8_2 & bh3_w8_3 & bh3_w8_4 & bh3_w8_5;
   Compressor_6_3_F800_uid6_uid43: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid43_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid43_Out0_copy44);
   Compressor_6_3_F800_uid6_bh3_uid43_Out0 <= Compressor_6_3_F800_uid6_bh3_uid43_Out0_copy44; -- output copy to hold a pipeline register if needed

   bh3_w8_14 <= Compressor_6_3_F800_uid6_bh3_uid43_Out0(0);
   bh3_w9_11 <= Compressor_6_3_F800_uid6_bh3_uid43_Out0(1);
   bh3_w10_10 <= Compressor_6_3_F800_uid6_bh3_uid43_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid45_In0 <= "" & bh3_w8_6 & bh3_w8_7 & bh3_w8_8 & bh3_w8_9;
   Compressor_14_3_F800_uid10_bh3_uid45_In1 <= "" & bh3_w9_0;
   Compressor_14_3_F800_uid10_uid45: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid45_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid45_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid45_Out0_copy46);
   Compressor_14_3_F800_uid10_bh3_uid45_Out0 <= Compressor_14_3_F800_uid10_bh3_uid45_Out0_copy46; -- output copy to hold a pipeline register if needed

   bh3_w8_15 <= Compressor_14_3_F800_uid10_bh3_uid45_Out0(0);
   bh3_w9_12 <= Compressor_14_3_F800_uid10_bh3_uid45_Out0(1);
   bh3_w10_11 <= Compressor_14_3_F800_uid10_bh3_uid45_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid47_In0 <= "" & bh3_w9_1 & bh3_w9_2 & bh3_w9_3 & bh3_w9_4 & bh3_w9_5 & bh3_w9_6;
   Compressor_6_3_F800_uid6_uid47: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid47_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid47_Out0_copy48);
   Compressor_6_3_F800_uid6_bh3_uid47_Out0 <= Compressor_6_3_F800_uid6_bh3_uid47_Out0_copy48; -- output copy to hold a pipeline register if needed

   bh3_w9_13 <= Compressor_6_3_F800_uid6_bh3_uid47_Out0(0);
   bh3_w10_12 <= Compressor_6_3_F800_uid6_bh3_uid47_Out0(1);
   bh3_w11_10 <= Compressor_6_3_F800_uid6_bh3_uid47_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid49_In0 <= "" & bh3_w9_7 & bh3_w9_8 & bh3_w9_9;
   Compressor_3_2_F800_uid16_uid49: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid49_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid49_Out0_copy50);
   Compressor_3_2_F800_uid16_bh3_uid49_Out0 <= Compressor_3_2_F800_uid16_bh3_uid49_Out0_copy50; -- output copy to hold a pipeline register if needed

   bh3_w9_14 <= Compressor_3_2_F800_uid16_bh3_uid49_Out0(0);
   bh3_w10_13 <= Compressor_3_2_F800_uid16_bh3_uid49_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid51_In0 <= "" & bh3_w10_0 & bh3_w10_1 & bh3_w10_2 & bh3_w10_3 & bh3_w10_4 & bh3_w10_5;
   Compressor_6_3_F800_uid6_uid51: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid51_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid51_Out0_copy52);
   Compressor_6_3_F800_uid6_bh3_uid51_Out0 <= Compressor_6_3_F800_uid6_bh3_uid51_Out0_copy52; -- output copy to hold a pipeline register if needed

   bh3_w10_14 <= Compressor_6_3_F800_uid6_bh3_uid51_Out0(0);
   bh3_w11_11 <= Compressor_6_3_F800_uid6_bh3_uid51_Out0(1);
   bh3_w12_10 <= Compressor_6_3_F800_uid6_bh3_uid51_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid53_In0 <= "" & bh3_w10_6 & bh3_w10_7 & bh3_w10_8 & bh3_w10_9;
   Compressor_14_3_F800_uid10_bh3_uid53_In1 <= "" & bh3_w11_0;
   Compressor_14_3_F800_uid10_uid53: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid53_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid53_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid53_Out0_copy54);
   Compressor_14_3_F800_uid10_bh3_uid53_Out0 <= Compressor_14_3_F800_uid10_bh3_uid53_Out0_copy54; -- output copy to hold a pipeline register if needed

   bh3_w10_15 <= Compressor_14_3_F800_uid10_bh3_uid53_Out0(0);
   bh3_w11_12 <= Compressor_14_3_F800_uid10_bh3_uid53_Out0(1);
   bh3_w12_11 <= Compressor_14_3_F800_uid10_bh3_uid53_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid55_In0 <= "" & bh3_w11_1 & bh3_w11_2 & bh3_w11_3 & bh3_w11_4 & bh3_w11_5 & bh3_w11_6;
   Compressor_6_3_F800_uid6_uid55: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid55_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid55_Out0_copy56);
   Compressor_6_3_F800_uid6_bh3_uid55_Out0 <= Compressor_6_3_F800_uid6_bh3_uid55_Out0_copy56; -- output copy to hold a pipeline register if needed

   bh3_w11_13 <= Compressor_6_3_F800_uid6_bh3_uid55_Out0(0);
   bh3_w12_12 <= Compressor_6_3_F800_uid6_bh3_uid55_Out0(1);
   bh3_w13_10 <= Compressor_6_3_F800_uid6_bh3_uid55_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid57_In0 <= "" & bh3_w11_7 & bh3_w11_8 & bh3_w11_9;
   Compressor_3_2_F800_uid16_uid57: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid57_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid57_Out0_copy58);
   Compressor_3_2_F800_uid16_bh3_uid57_Out0 <= Compressor_3_2_F800_uid16_bh3_uid57_Out0_copy58; -- output copy to hold a pipeline register if needed

   bh3_w11_14 <= Compressor_3_2_F800_uid16_bh3_uid57_Out0(0);
   bh3_w12_13 <= Compressor_3_2_F800_uid16_bh3_uid57_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid59_In0 <= "" & bh3_w12_0 & bh3_w12_1 & bh3_w12_2 & bh3_w12_3 & bh3_w12_4 & bh3_w12_5;
   Compressor_6_3_F800_uid6_uid59: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid59_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid59_Out0_copy60);
   Compressor_6_3_F800_uid6_bh3_uid59_Out0 <= Compressor_6_3_F800_uid6_bh3_uid59_Out0_copy60; -- output copy to hold a pipeline register if needed

   bh3_w12_14 <= Compressor_6_3_F800_uid6_bh3_uid59_Out0(0);
   bh3_w13_11 <= Compressor_6_3_F800_uid6_bh3_uid59_Out0(1);
   bh3_w14_10 <= Compressor_6_3_F800_uid6_bh3_uid59_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid61_In0 <= "" & bh3_w12_6 & bh3_w12_7 & bh3_w12_8 & bh3_w12_9;
   Compressor_14_3_F800_uid10_bh3_uid61_In1 <= "" & bh3_w13_0;
   Compressor_14_3_F800_uid10_uid61: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid61_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid61_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid61_Out0_copy62);
   Compressor_14_3_F800_uid10_bh3_uid61_Out0 <= Compressor_14_3_F800_uid10_bh3_uid61_Out0_copy62; -- output copy to hold a pipeline register if needed

   bh3_w12_15 <= Compressor_14_3_F800_uid10_bh3_uid61_Out0(0);
   bh3_w13_12 <= Compressor_14_3_F800_uid10_bh3_uid61_Out0(1);
   bh3_w14_11 <= Compressor_14_3_F800_uid10_bh3_uid61_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid63_In0 <= "" & bh3_w13_1 & bh3_w13_2 & bh3_w13_3 & bh3_w13_4 & bh3_w13_5 & bh3_w13_6;
   Compressor_6_3_F800_uid6_uid63: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid63_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid63_Out0_copy64);
   Compressor_6_3_F800_uid6_bh3_uid63_Out0 <= Compressor_6_3_F800_uid6_bh3_uid63_Out0_copy64; -- output copy to hold a pipeline register if needed

   bh3_w13_13 <= Compressor_6_3_F800_uid6_bh3_uid63_Out0(0);
   bh3_w14_12 <= Compressor_6_3_F800_uid6_bh3_uid63_Out0(1);
   bh3_w15_10 <= Compressor_6_3_F800_uid6_bh3_uid63_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid65_In0 <= "" & bh3_w13_7 & bh3_w13_8 & bh3_w13_9;
   Compressor_3_2_F800_uid16_uid65: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid65_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid65_Out0_copy66);
   Compressor_3_2_F800_uid16_bh3_uid65_Out0 <= Compressor_3_2_F800_uid16_bh3_uid65_Out0_copy66; -- output copy to hold a pipeline register if needed

   bh3_w13_14 <= Compressor_3_2_F800_uid16_bh3_uid65_Out0(0);
   bh3_w14_13 <= Compressor_3_2_F800_uid16_bh3_uid65_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid67_In0 <= "" & bh3_w14_0 & bh3_w14_1 & bh3_w14_2 & bh3_w14_3 & bh3_w14_4 & bh3_w14_5;
   Compressor_6_3_F800_uid6_uid67: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid67_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid67_Out0_copy68);
   Compressor_6_3_F800_uid6_bh3_uid67_Out0 <= Compressor_6_3_F800_uid6_bh3_uid67_Out0_copy68; -- output copy to hold a pipeline register if needed

   bh3_w14_14 <= Compressor_6_3_F800_uid6_bh3_uid67_Out0(0);
   bh3_w15_11 <= Compressor_6_3_F800_uid6_bh3_uid67_Out0(1);
   bh3_w16_10 <= Compressor_6_3_F800_uid6_bh3_uid67_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid69_In0 <= "" & bh3_w14_6 & bh3_w14_7 & bh3_w14_8 & bh3_w14_9;
   Compressor_14_3_F800_uid10_bh3_uid69_In1 <= "" & bh3_w15_0;
   Compressor_14_3_F800_uid10_uid69: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid69_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid69_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid69_Out0_copy70);
   Compressor_14_3_F800_uid10_bh3_uid69_Out0 <= Compressor_14_3_F800_uid10_bh3_uid69_Out0_copy70; -- output copy to hold a pipeline register if needed

   bh3_w14_15 <= Compressor_14_3_F800_uid10_bh3_uid69_Out0(0);
   bh3_w15_12 <= Compressor_14_3_F800_uid10_bh3_uid69_Out0(1);
   bh3_w16_11 <= Compressor_14_3_F800_uid10_bh3_uid69_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid71_In0 <= "" & bh3_w15_1 & bh3_w15_2 & bh3_w15_3 & bh3_w15_4 & bh3_w15_5 & bh3_w15_6;
   Compressor_6_3_F800_uid6_uid71: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid71_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid71_Out0_copy72);
   Compressor_6_3_F800_uid6_bh3_uid71_Out0 <= Compressor_6_3_F800_uid6_bh3_uid71_Out0_copy72; -- output copy to hold a pipeline register if needed

   bh3_w15_13 <= Compressor_6_3_F800_uid6_bh3_uid71_Out0(0);
   bh3_w16_12 <= Compressor_6_3_F800_uid6_bh3_uid71_Out0(1);
   bh3_w17_10 <= Compressor_6_3_F800_uid6_bh3_uid71_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid73_In0 <= "" & bh3_w15_7 & bh3_w15_8 & bh3_w15_9;
   Compressor_3_2_F800_uid16_uid73: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid73_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid73_Out0_copy74);
   Compressor_3_2_F800_uid16_bh3_uid73_Out0 <= Compressor_3_2_F800_uid16_bh3_uid73_Out0_copy74; -- output copy to hold a pipeline register if needed

   bh3_w15_14 <= Compressor_3_2_F800_uid16_bh3_uid73_Out0(0);
   bh3_w16_13 <= Compressor_3_2_F800_uid16_bh3_uid73_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid75_In0 <= "" & bh3_w16_0 & bh3_w16_1 & bh3_w16_2 & bh3_w16_3 & bh3_w16_4 & bh3_w16_5;
   Compressor_6_3_F800_uid6_uid75: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid75_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid75_Out0_copy76);
   Compressor_6_3_F800_uid6_bh3_uid75_Out0 <= Compressor_6_3_F800_uid6_bh3_uid75_Out0_copy76; -- output copy to hold a pipeline register if needed

   bh3_w16_14 <= Compressor_6_3_F800_uid6_bh3_uid75_Out0(0);
   bh3_w17_11 <= Compressor_6_3_F800_uid6_bh3_uid75_Out0(1);
   bh3_w18_10 <= Compressor_6_3_F800_uid6_bh3_uid75_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid77_In0 <= "" & bh3_w16_6 & bh3_w16_7 & bh3_w16_8 & bh3_w16_9;
   Compressor_14_3_F800_uid10_bh3_uid77_In1 <= "" & bh3_w17_0;
   Compressor_14_3_F800_uid10_uid77: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid77_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid77_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid77_Out0_copy78);
   Compressor_14_3_F800_uid10_bh3_uid77_Out0 <= Compressor_14_3_F800_uid10_bh3_uid77_Out0_copy78; -- output copy to hold a pipeline register if needed

   bh3_w16_15 <= Compressor_14_3_F800_uid10_bh3_uid77_Out0(0);
   bh3_w17_12 <= Compressor_14_3_F800_uid10_bh3_uid77_Out0(1);
   bh3_w18_11 <= Compressor_14_3_F800_uid10_bh3_uid77_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid79_In0 <= "" & bh3_w17_1 & bh3_w17_2 & bh3_w17_3 & bh3_w17_4 & bh3_w17_5 & bh3_w17_6;
   Compressor_6_3_F800_uid6_uid79: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid79_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid79_Out0_copy80);
   Compressor_6_3_F800_uid6_bh3_uid79_Out0 <= Compressor_6_3_F800_uid6_bh3_uid79_Out0_copy80; -- output copy to hold a pipeline register if needed

   bh3_w17_13 <= Compressor_6_3_F800_uid6_bh3_uid79_Out0(0);
   bh3_w18_12 <= Compressor_6_3_F800_uid6_bh3_uid79_Out0(1);
   bh3_w19_10 <= Compressor_6_3_F800_uid6_bh3_uid79_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid81_In0 <= "" & bh3_w17_7 & bh3_w17_8 & bh3_w17_9;
   Compressor_3_2_F800_uid16_uid81: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid81_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid81_Out0_copy82);
   Compressor_3_2_F800_uid16_bh3_uid81_Out0 <= Compressor_3_2_F800_uid16_bh3_uid81_Out0_copy82; -- output copy to hold a pipeline register if needed

   bh3_w17_14 <= Compressor_3_2_F800_uid16_bh3_uid81_Out0(0);
   bh3_w18_13 <= Compressor_3_2_F800_uid16_bh3_uid81_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid83_In0 <= "" & bh3_w18_0 & bh3_w18_1 & bh3_w18_2 & bh3_w18_3 & bh3_w18_4 & bh3_w18_5;
   Compressor_6_3_F800_uid6_uid83: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid83_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid83_Out0_copy84);
   Compressor_6_3_F800_uid6_bh3_uid83_Out0 <= Compressor_6_3_F800_uid6_bh3_uid83_Out0_copy84; -- output copy to hold a pipeline register if needed

   bh3_w18_14 <= Compressor_6_3_F800_uid6_bh3_uid83_Out0(0);
   bh3_w19_11 <= Compressor_6_3_F800_uid6_bh3_uid83_Out0(1);
   bh3_w20_0 <= Compressor_6_3_F800_uid6_bh3_uid83_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid85_In0 <= "" & bh3_w18_6 & bh3_w18_7 & bh3_w18_8 & bh3_w18_9;
   Compressor_14_3_F800_uid10_bh3_uid85_In1 <= "" & bh3_w19_0;
   Compressor_14_3_F800_uid10_uid85: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid85_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid85_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid85_Out0_copy86);
   Compressor_14_3_F800_uid10_bh3_uid85_Out0 <= Compressor_14_3_F800_uid10_bh3_uid85_Out0_copy86; -- output copy to hold a pipeline register if needed

   bh3_w18_15 <= Compressor_14_3_F800_uid10_bh3_uid85_Out0(0);
   bh3_w19_12 <= Compressor_14_3_F800_uid10_bh3_uid85_Out0(1);
   bh3_w20_1 <= Compressor_14_3_F800_uid10_bh3_uid85_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid87_In0 <= "" & bh3_w19_1 & bh3_w19_2 & bh3_w19_3 & bh3_w19_4 & bh3_w19_5 & bh3_w19_6;
   Compressor_6_3_F800_uid6_uid87: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid87_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid87_Out0_copy88);
   Compressor_6_3_F800_uid6_bh3_uid87_Out0 <= Compressor_6_3_F800_uid6_bh3_uid87_Out0_copy88; -- output copy to hold a pipeline register if needed

   bh3_w19_13 <= Compressor_6_3_F800_uid6_bh3_uid87_Out0(0);
   bh3_w20_2 <= Compressor_6_3_F800_uid6_bh3_uid87_Out0(1);
   bh3_w21_0 <= Compressor_6_3_F800_uid6_bh3_uid87_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid89_In0 <= "" & bh3_w19_7 & bh3_w19_8 & bh3_w19_9;
   Compressor_3_2_F800_uid16_uid89: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid89_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid89_Out0_copy90);
   Compressor_3_2_F800_uid16_bh3_uid89_Out0 <= Compressor_3_2_F800_uid16_bh3_uid89_Out0_copy90; -- output copy to hold a pipeline register if needed

   bh3_w19_14 <= Compressor_3_2_F800_uid16_bh3_uid89_Out0(0);
   bh3_w20_3 <= Compressor_3_2_F800_uid16_bh3_uid89_Out0(1);

   Compressor_14_3_F800_uid10_bh3_uid91_In0 <= "" & bh3_w0_11 & bh3_w0_10 & "0" & "0";
   Compressor_14_3_F800_uid10_bh3_uid91_In1 <= "" & bh3_w1_13;
   Compressor_14_3_F800_uid10_uid91: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid91_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid91_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92);
   Compressor_14_3_F800_uid10_bh3_uid91_Out0 <= Compressor_14_3_F800_uid10_bh3_uid91_Out0_copy92_d1; -- output copy to hold a pipeline register if needed

   bh3_w0_12 <= Compressor_14_3_F800_uid10_bh3_uid91_Out0(0);
   bh3_w1_14 <= Compressor_14_3_F800_uid10_bh3_uid91_Out0(1);
   bh3_w2_16 <= Compressor_14_3_F800_uid10_bh3_uid91_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid93_In0 <= "" & bh3_w1_12 & bh3_w1_11 & bh3_w1_10;
   Compressor_3_2_F800_uid16_uid93: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid93_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94);
   Compressor_3_2_F800_uid16_bh3_uid93_Out0 <= Compressor_3_2_F800_uid16_bh3_uid93_Out0_copy94_d1; -- output copy to hold a pipeline register if needed

   bh3_w1_15 <= Compressor_3_2_F800_uid16_bh3_uid93_Out0(0);
   bh3_w2_17 <= Compressor_3_2_F800_uid16_bh3_uid93_Out0(1);

   Compressor_6_3_F800_uid6_bh3_uid95_In0 <= "" & bh3_w2_15 & bh3_w2_14 & bh3_w2_13 & bh3_w2_12 & bh3_w2_11 & bh3_w2_10;
   Compressor_6_3_F800_uid6_uid95: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid95_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96);
   Compressor_6_3_F800_uid6_bh3_uid95_Out0 <= Compressor_6_3_F800_uid6_bh3_uid95_Out0_copy96_d1; -- output copy to hold a pipeline register if needed

   bh3_w2_18 <= Compressor_6_3_F800_uid6_bh3_uid95_Out0(0);
   bh3_w3_15 <= Compressor_6_3_F800_uid6_bh3_uid95_Out0(1);
   bh3_w4_16 <= Compressor_6_3_F800_uid6_bh3_uid95_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid99_In0 <= "" & bh3_w3_14 & bh3_w3_13 & bh3_w3_12 & bh3_w3_11 & bh3_w3_10;
   Compressor_5_3_F800_uid98_uid99: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid99_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100);
   Compressor_5_3_F800_uid98_bh3_uid99_Out0 <= Compressor_5_3_F800_uid98_bh3_uid99_Out0_copy100_d1; -- output copy to hold a pipeline register if needed

   bh3_w3_16 <= Compressor_5_3_F800_uid98_bh3_uid99_Out0(0);
   bh3_w4_17 <= Compressor_5_3_F800_uid98_bh3_uid99_Out0(1);
   bh3_w5_15 <= Compressor_5_3_F800_uid98_bh3_uid99_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid101_In0 <= "" & bh3_w4_15 & bh3_w4_14 & bh3_w4_13 & bh3_w4_12 & bh3_w4_11 & bh3_w4_10;
   Compressor_6_3_F800_uid6_uid101: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid101_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102);
   Compressor_6_3_F800_uid6_bh3_uid101_Out0 <= Compressor_6_3_F800_uid6_bh3_uid101_Out0_copy102_d1; -- output copy to hold a pipeline register if needed

   bh3_w4_18 <= Compressor_6_3_F800_uid6_bh3_uid101_Out0(0);
   bh3_w5_16 <= Compressor_6_3_F800_uid6_bh3_uid101_Out0(1);
   bh3_w6_16 <= Compressor_6_3_F800_uid6_bh3_uid101_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid103_In0 <= "" & bh3_w5_14 & bh3_w5_13 & bh3_w5_12 & bh3_w5_11 & bh3_w5_10;
   Compressor_5_3_F800_uid98_uid103: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid103_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104);
   Compressor_5_3_F800_uid98_bh3_uid103_Out0 <= Compressor_5_3_F800_uid98_bh3_uid103_Out0_copy104_d1; -- output copy to hold a pipeline register if needed

   bh3_w5_17 <= Compressor_5_3_F800_uid98_bh3_uid103_Out0(0);
   bh3_w6_17 <= Compressor_5_3_F800_uid98_bh3_uid103_Out0(1);
   bh3_w7_15 <= Compressor_5_3_F800_uid98_bh3_uid103_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid105_In0 <= "" & bh3_w6_15 & bh3_w6_14 & bh3_w6_13 & bh3_w6_12 & bh3_w6_11 & bh3_w6_10;
   Compressor_6_3_F800_uid6_uid105: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid105_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106);
   Compressor_6_3_F800_uid6_bh3_uid105_Out0 <= Compressor_6_3_F800_uid6_bh3_uid105_Out0_copy106_d1; -- output copy to hold a pipeline register if needed

   bh3_w6_18 <= Compressor_6_3_F800_uid6_bh3_uid105_Out0(0);
   bh3_w7_16 <= Compressor_6_3_F800_uid6_bh3_uid105_Out0(1);
   bh3_w8_16 <= Compressor_6_3_F800_uid6_bh3_uid105_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid107_In0 <= "" & bh3_w7_14 & bh3_w7_13 & bh3_w7_12 & bh3_w7_11 & bh3_w7_10;
   Compressor_5_3_F800_uid98_uid107: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid107_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108);
   Compressor_5_3_F800_uid98_bh3_uid107_Out0 <= Compressor_5_3_F800_uid98_bh3_uid107_Out0_copy108_d1; -- output copy to hold a pipeline register if needed

   bh3_w7_17 <= Compressor_5_3_F800_uid98_bh3_uid107_Out0(0);
   bh3_w8_17 <= Compressor_5_3_F800_uid98_bh3_uid107_Out0(1);
   bh3_w9_15 <= Compressor_5_3_F800_uid98_bh3_uid107_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid109_In0 <= "" & bh3_w8_15 & bh3_w8_14 & bh3_w8_13 & bh3_w8_12 & bh3_w8_11 & bh3_w8_10;
   Compressor_6_3_F800_uid6_uid109: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid109_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110);
   Compressor_6_3_F800_uid6_bh3_uid109_Out0 <= Compressor_6_3_F800_uid6_bh3_uid109_Out0_copy110_d1; -- output copy to hold a pipeline register if needed

   bh3_w8_18 <= Compressor_6_3_F800_uid6_bh3_uid109_Out0(0);
   bh3_w9_16 <= Compressor_6_3_F800_uid6_bh3_uid109_Out0(1);
   bh3_w10_16 <= Compressor_6_3_F800_uid6_bh3_uid109_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid111_In0 <= "" & bh3_w9_14 & bh3_w9_13 & bh3_w9_12 & bh3_w9_11 & bh3_w9_10;
   Compressor_5_3_F800_uid98_uid111: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid111_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112);
   Compressor_5_3_F800_uid98_bh3_uid111_Out0 <= Compressor_5_3_F800_uid98_bh3_uid111_Out0_copy112_d1; -- output copy to hold a pipeline register if needed

   bh3_w9_17 <= Compressor_5_3_F800_uid98_bh3_uid111_Out0(0);
   bh3_w10_17 <= Compressor_5_3_F800_uid98_bh3_uid111_Out0(1);
   bh3_w11_15 <= Compressor_5_3_F800_uid98_bh3_uid111_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid113_In0 <= "" & bh3_w10_15 & bh3_w10_14 & bh3_w10_13 & bh3_w10_12 & bh3_w10_11 & bh3_w10_10;
   Compressor_6_3_F800_uid6_uid113: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid113_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114);
   Compressor_6_3_F800_uid6_bh3_uid113_Out0 <= Compressor_6_3_F800_uid6_bh3_uid113_Out0_copy114_d1; -- output copy to hold a pipeline register if needed

   bh3_w10_18 <= Compressor_6_3_F800_uid6_bh3_uid113_Out0(0);
   bh3_w11_16 <= Compressor_6_3_F800_uid6_bh3_uid113_Out0(1);
   bh3_w12_16 <= Compressor_6_3_F800_uid6_bh3_uid113_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid115_In0 <= "" & bh3_w11_14 & bh3_w11_13 & bh3_w11_12 & bh3_w11_11 & bh3_w11_10;
   Compressor_5_3_F800_uid98_uid115: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid115_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116);
   Compressor_5_3_F800_uid98_bh3_uid115_Out0 <= Compressor_5_3_F800_uid98_bh3_uid115_Out0_copy116_d1; -- output copy to hold a pipeline register if needed

   bh3_w11_17 <= Compressor_5_3_F800_uid98_bh3_uid115_Out0(0);
   bh3_w12_17 <= Compressor_5_3_F800_uid98_bh3_uid115_Out0(1);
   bh3_w13_15 <= Compressor_5_3_F800_uid98_bh3_uid115_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid117_In0 <= "" & bh3_w12_15 & bh3_w12_14 & bh3_w12_13 & bh3_w12_12 & bh3_w12_11 & bh3_w12_10;
   Compressor_6_3_F800_uid6_uid117: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid117_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118);
   Compressor_6_3_F800_uid6_bh3_uid117_Out0 <= Compressor_6_3_F800_uid6_bh3_uid117_Out0_copy118_d1; -- output copy to hold a pipeline register if needed

   bh3_w12_18 <= Compressor_6_3_F800_uid6_bh3_uid117_Out0(0);
   bh3_w13_16 <= Compressor_6_3_F800_uid6_bh3_uid117_Out0(1);
   bh3_w14_16 <= Compressor_6_3_F800_uid6_bh3_uid117_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid119_In0 <= "" & bh3_w13_14 & bh3_w13_13 & bh3_w13_12 & bh3_w13_11 & bh3_w13_10;
   Compressor_5_3_F800_uid98_uid119: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid119_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120);
   Compressor_5_3_F800_uid98_bh3_uid119_Out0 <= Compressor_5_3_F800_uid98_bh3_uid119_Out0_copy120_d1; -- output copy to hold a pipeline register if needed

   bh3_w13_17 <= Compressor_5_3_F800_uid98_bh3_uid119_Out0(0);
   bh3_w14_17 <= Compressor_5_3_F800_uid98_bh3_uid119_Out0(1);
   bh3_w15_15 <= Compressor_5_3_F800_uid98_bh3_uid119_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid121_In0 <= "" & bh3_w14_15 & bh3_w14_14 & bh3_w14_13 & bh3_w14_12 & bh3_w14_11 & bh3_w14_10;
   Compressor_6_3_F800_uid6_uid121: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid121_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122);
   Compressor_6_3_F800_uid6_bh3_uid121_Out0 <= Compressor_6_3_F800_uid6_bh3_uid121_Out0_copy122_d1; -- output copy to hold a pipeline register if needed

   bh3_w14_18 <= Compressor_6_3_F800_uid6_bh3_uid121_Out0(0);
   bh3_w15_16 <= Compressor_6_3_F800_uid6_bh3_uid121_Out0(1);
   bh3_w16_16 <= Compressor_6_3_F800_uid6_bh3_uid121_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid123_In0 <= "" & bh3_w15_14 & bh3_w15_13 & bh3_w15_12 & bh3_w15_11 & bh3_w15_10;
   Compressor_5_3_F800_uid98_uid123: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid123_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124);
   Compressor_5_3_F800_uid98_bh3_uid123_Out0 <= Compressor_5_3_F800_uid98_bh3_uid123_Out0_copy124_d1; -- output copy to hold a pipeline register if needed

   bh3_w15_17 <= Compressor_5_3_F800_uid98_bh3_uid123_Out0(0);
   bh3_w16_17 <= Compressor_5_3_F800_uid98_bh3_uid123_Out0(1);
   bh3_w17_15 <= Compressor_5_3_F800_uid98_bh3_uid123_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid125_In0 <= "" & bh3_w16_15 & bh3_w16_14 & bh3_w16_13 & bh3_w16_12 & bh3_w16_11 & bh3_w16_10;
   Compressor_6_3_F800_uid6_uid125: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid125_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126);
   Compressor_6_3_F800_uid6_bh3_uid125_Out0 <= Compressor_6_3_F800_uid6_bh3_uid125_Out0_copy126_d1; -- output copy to hold a pipeline register if needed

   bh3_w16_18 <= Compressor_6_3_F800_uid6_bh3_uid125_Out0(0);
   bh3_w17_16 <= Compressor_6_3_F800_uid6_bh3_uid125_Out0(1);
   bh3_w18_16 <= Compressor_6_3_F800_uid6_bh3_uid125_Out0(2);

   Compressor_5_3_F800_uid98_bh3_uid127_In0 <= "" & bh3_w17_14 & bh3_w17_13 & bh3_w17_12 & bh3_w17_11 & bh3_w17_10;
   Compressor_5_3_F800_uid98_uid127: Compressor_5_3_F800_uid98
      port map ( X0 => Compressor_5_3_F800_uid98_bh3_uid127_In0,
                 R => Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128);
   Compressor_5_3_F800_uid98_bh3_uid127_Out0 <= Compressor_5_3_F800_uid98_bh3_uid127_Out0_copy128_d1; -- output copy to hold a pipeline register if needed

   bh3_w17_17 <= Compressor_5_3_F800_uid98_bh3_uid127_Out0(0);
   bh3_w18_17 <= Compressor_5_3_F800_uid98_bh3_uid127_Out0(1);
   bh3_w19_15 <= Compressor_5_3_F800_uid98_bh3_uid127_Out0(2);

   Compressor_6_3_F800_uid6_bh3_uid129_In0 <= "" & bh3_w18_15 & bh3_w18_14 & bh3_w18_13 & bh3_w18_12 & bh3_w18_11 & bh3_w18_10;
   Compressor_6_3_F800_uid6_uid129: Compressor_6_3_F800_uid6
      port map ( X0 => Compressor_6_3_F800_uid6_bh3_uid129_In0,
                 R => Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130);
   Compressor_6_3_F800_uid6_bh3_uid129_Out0 <= Compressor_6_3_F800_uid6_bh3_uid129_Out0_copy130_d1; -- output copy to hold a pipeline register if needed

   bh3_w18_18 <= Compressor_6_3_F800_uid6_bh3_uid129_Out0(0);
   bh3_w19_16 <= Compressor_6_3_F800_uid6_bh3_uid129_Out0(1);
   bh3_w20_4 <= Compressor_6_3_F800_uid6_bh3_uid129_Out0(2);

   Compressor_14_3_F800_uid10_bh3_uid131_In0 <= "" & bh3_w19_14 & bh3_w19_13 & bh3_w19_12 & bh3_w19_11;
   Compressor_14_3_F800_uid10_bh3_uid131_In1 <= "" & bh3_w20_3;
   Compressor_14_3_F800_uid10_uid131: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid131_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid131_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132);
   Compressor_14_3_F800_uid10_bh3_uid131_Out0 <= Compressor_14_3_F800_uid10_bh3_uid131_Out0_copy132_d1; -- output copy to hold a pipeline register if needed

   bh3_w19_17 <= Compressor_14_3_F800_uid10_bh3_uid131_Out0(0);
   bh3_w20_5 <= Compressor_14_3_F800_uid10_bh3_uid131_Out0(1);
   bh3_w21_1 <= Compressor_14_3_F800_uid10_bh3_uid131_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid133_In0 <= "" & bh3_w20_2 & bh3_w20_1 & bh3_w20_0;
   Compressor_3_2_F800_uid16_uid133: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid133_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134);
   Compressor_3_2_F800_uid16_bh3_uid133_Out0 <= Compressor_3_2_F800_uid16_bh3_uid133_Out0_copy134_d1; -- output copy to hold a pipeline register if needed

   bh3_w20_6 <= Compressor_3_2_F800_uid16_bh3_uid133_Out0(0);
   bh3_w21_2 <= Compressor_3_2_F800_uid16_bh3_uid133_Out0(1);

   Compressor_23_3_F800_uid136_bh3_uid137_In0 <= "" & bh3_w0_12 & "0" & "0";
   Compressor_23_3_F800_uid136_bh3_uid137_In1 <= "" & bh3_w1_15 & bh3_w1_14;
   Compressor_23_3_F800_uid136_uid137: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid137_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid137_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid137_Out0_copy138);
   Compressor_23_3_F800_uid136_bh3_uid137_Out0 <= Compressor_23_3_F800_uid136_bh3_uid137_Out0_copy138; -- output copy to hold a pipeline register if needed

   bh3_w0_13 <= Compressor_23_3_F800_uid136_bh3_uid137_Out0(0);
   bh3_w1_16 <= Compressor_23_3_F800_uid136_bh3_uid137_Out0(1);
   bh3_w2_19 <= Compressor_23_3_F800_uid136_bh3_uid137_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid139_In0 <= "" & bh3_w2_18 & bh3_w2_17 & bh3_w2_16;
   Compressor_23_3_F800_uid136_bh3_uid139_In1 <= "" & bh3_w3_16 & bh3_w3_15;
   Compressor_23_3_F800_uid136_uid139: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid139_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid139_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid139_Out0_copy140);
   Compressor_23_3_F800_uid136_bh3_uid139_Out0 <= Compressor_23_3_F800_uid136_bh3_uid139_Out0_copy140; -- output copy to hold a pipeline register if needed

   bh3_w2_20 <= Compressor_23_3_F800_uid136_bh3_uid139_Out0(0);
   bh3_w3_17 <= Compressor_23_3_F800_uid136_bh3_uid139_Out0(1);
   bh3_w4_19 <= Compressor_23_3_F800_uid136_bh3_uid139_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid141_In0 <= "" & bh3_w4_18 & bh3_w4_17 & bh3_w4_16;
   Compressor_23_3_F800_uid136_bh3_uid141_In1 <= "" & bh3_w5_17 & bh3_w5_16;
   Compressor_23_3_F800_uid136_uid141: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid141_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid141_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid141_Out0_copy142);
   Compressor_23_3_F800_uid136_bh3_uid141_Out0 <= Compressor_23_3_F800_uid136_bh3_uid141_Out0_copy142; -- output copy to hold a pipeline register if needed

   bh3_w4_20 <= Compressor_23_3_F800_uid136_bh3_uid141_Out0(0);
   bh3_w5_18 <= Compressor_23_3_F800_uid136_bh3_uid141_Out0(1);
   bh3_w6_19 <= Compressor_23_3_F800_uid136_bh3_uid141_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid143_In0 <= "" & bh3_w6_18 & bh3_w6_17 & bh3_w6_16;
   Compressor_23_3_F800_uid136_bh3_uid143_In1 <= "" & bh3_w7_17 & bh3_w7_16;
   Compressor_23_3_F800_uid136_uid143: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid143_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid143_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid143_Out0_copy144);
   Compressor_23_3_F800_uid136_bh3_uid143_Out0 <= Compressor_23_3_F800_uid136_bh3_uid143_Out0_copy144; -- output copy to hold a pipeline register if needed

   bh3_w6_20 <= Compressor_23_3_F800_uid136_bh3_uid143_Out0(0);
   bh3_w7_18 <= Compressor_23_3_F800_uid136_bh3_uid143_Out0(1);
   bh3_w8_19 <= Compressor_23_3_F800_uid136_bh3_uid143_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid145_In0 <= "" & bh3_w8_18 & bh3_w8_17 & bh3_w8_16;
   Compressor_23_3_F800_uid136_bh3_uid145_In1 <= "" & bh3_w9_17 & bh3_w9_16;
   Compressor_23_3_F800_uid136_uid145: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid145_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid145_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid145_Out0_copy146);
   Compressor_23_3_F800_uid136_bh3_uid145_Out0 <= Compressor_23_3_F800_uid136_bh3_uid145_Out0_copy146; -- output copy to hold a pipeline register if needed

   bh3_w8_20 <= Compressor_23_3_F800_uid136_bh3_uid145_Out0(0);
   bh3_w9_18 <= Compressor_23_3_F800_uid136_bh3_uid145_Out0(1);
   bh3_w10_19 <= Compressor_23_3_F800_uid136_bh3_uid145_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid147_In0 <= "" & bh3_w10_18 & bh3_w10_17 & bh3_w10_16;
   Compressor_23_3_F800_uid136_bh3_uid147_In1 <= "" & bh3_w11_17 & bh3_w11_16;
   Compressor_23_3_F800_uid136_uid147: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid147_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid147_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid147_Out0_copy148);
   Compressor_23_3_F800_uid136_bh3_uid147_Out0 <= Compressor_23_3_F800_uid136_bh3_uid147_Out0_copy148; -- output copy to hold a pipeline register if needed

   bh3_w10_20 <= Compressor_23_3_F800_uid136_bh3_uid147_Out0(0);
   bh3_w11_18 <= Compressor_23_3_F800_uid136_bh3_uid147_Out0(1);
   bh3_w12_19 <= Compressor_23_3_F800_uid136_bh3_uid147_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid149_In0 <= "" & bh3_w12_18 & bh3_w12_17 & bh3_w12_16;
   Compressor_23_3_F800_uid136_bh3_uid149_In1 <= "" & bh3_w13_17 & bh3_w13_16;
   Compressor_23_3_F800_uid136_uid149: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid149_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid149_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid149_Out0_copy150);
   Compressor_23_3_F800_uid136_bh3_uid149_Out0 <= Compressor_23_3_F800_uid136_bh3_uid149_Out0_copy150; -- output copy to hold a pipeline register if needed

   bh3_w12_20 <= Compressor_23_3_F800_uid136_bh3_uid149_Out0(0);
   bh3_w13_18 <= Compressor_23_3_F800_uid136_bh3_uid149_Out0(1);
   bh3_w14_19 <= Compressor_23_3_F800_uid136_bh3_uid149_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid151_In0 <= "" & bh3_w14_18 & bh3_w14_17 & bh3_w14_16;
   Compressor_23_3_F800_uid136_bh3_uid151_In1 <= "" & bh3_w15_17 & bh3_w15_16;
   Compressor_23_3_F800_uid136_uid151: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid151_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid151_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid151_Out0_copy152);
   Compressor_23_3_F800_uid136_bh3_uid151_Out0 <= Compressor_23_3_F800_uid136_bh3_uid151_Out0_copy152; -- output copy to hold a pipeline register if needed

   bh3_w14_20 <= Compressor_23_3_F800_uid136_bh3_uid151_Out0(0);
   bh3_w15_18 <= Compressor_23_3_F800_uid136_bh3_uid151_Out0(1);
   bh3_w16_19 <= Compressor_23_3_F800_uid136_bh3_uid151_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid153_In0 <= "" & bh3_w16_18 & bh3_w16_17 & bh3_w16_16;
   Compressor_23_3_F800_uid136_bh3_uid153_In1 <= "" & bh3_w17_17 & bh3_w17_16;
   Compressor_23_3_F800_uid136_uid153: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid153_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid153_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid153_Out0_copy154);
   Compressor_23_3_F800_uid136_bh3_uid153_Out0 <= Compressor_23_3_F800_uid136_bh3_uid153_Out0_copy154; -- output copy to hold a pipeline register if needed

   bh3_w16_20 <= Compressor_23_3_F800_uid136_bh3_uid153_Out0(0);
   bh3_w17_18 <= Compressor_23_3_F800_uid136_bh3_uid153_Out0(1);
   bh3_w18_19 <= Compressor_23_3_F800_uid136_bh3_uid153_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid155_In0 <= "" & bh3_w18_18 & bh3_w18_17 & bh3_w18_16;
   Compressor_3_2_F800_uid16_uid155: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid155_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid155_Out0_copy156);
   Compressor_3_2_F800_uid16_bh3_uid155_Out0 <= Compressor_3_2_F800_uid16_bh3_uid155_Out0_copy156; -- output copy to hold a pipeline register if needed

   bh3_w18_20 <= Compressor_3_2_F800_uid16_bh3_uid155_Out0(0);
   bh3_w19_18 <= Compressor_3_2_F800_uid16_bh3_uid155_Out0(1);

   Compressor_14_3_F800_uid10_bh3_uid157_In0 <= "" & bh3_w19_10_d1 & bh3_w19_17 & bh3_w19_16 & bh3_w19_15;
   Compressor_14_3_F800_uid10_bh3_uid157_In1 <= "" & "0";
   Compressor_14_3_F800_uid10_uid157: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid157_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid157_In1_d1,
                 R => Compressor_14_3_F800_uid10_bh3_uid157_Out0_copy158);
   Compressor_14_3_F800_uid10_bh3_uid157_Out0 <= Compressor_14_3_F800_uid10_bh3_uid157_Out0_copy158; -- output copy to hold a pipeline register if needed

   bh3_w19_19 <= Compressor_14_3_F800_uid10_bh3_uid157_Out0(0);
   bh3_w20_7 <= Compressor_14_3_F800_uid10_bh3_uid157_Out0(1);
   bh3_w21_3 <= Compressor_14_3_F800_uid10_bh3_uid157_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid159_In0 <= "" & bh3_w20_6 & bh3_w20_5 & bh3_w20_4;
   Compressor_3_2_F800_uid16_uid159: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid159_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid159_Out0_copy160);
   Compressor_3_2_F800_uid16_bh3_uid159_Out0 <= Compressor_3_2_F800_uid16_bh3_uid159_Out0_copy160; -- output copy to hold a pipeline register if needed

   bh3_w20_8 <= Compressor_3_2_F800_uid16_bh3_uid159_Out0(0);
   bh3_w21_4 <= Compressor_3_2_F800_uid16_bh3_uid159_Out0(1);

   Compressor_3_2_F800_uid16_bh3_uid161_In0 <= "" & bh3_w21_0_d1 & bh3_w21_2 & bh3_w21_1;
   Compressor_3_2_F800_uid16_uid161: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid161_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid161_Out0_copy162);
   Compressor_3_2_F800_uid16_bh3_uid161_Out0 <= Compressor_3_2_F800_uid16_bh3_uid161_Out0_copy162; -- output copy to hold a pipeline register if needed

   bh3_w21_5 <= Compressor_3_2_F800_uid16_bh3_uid161_Out0(0);
   bh3_w22_0 <= Compressor_3_2_F800_uid16_bh3_uid161_Out0(1);

   Compressor_14_3_F800_uid10_bh3_uid163_In0 <= "" & bh3_w2_20 & bh3_w2_19 & "0" & "0";
   Compressor_14_3_F800_uid10_bh3_uid163_In1 <= "" & bh3_w3_17;
   Compressor_14_3_F800_uid10_uid163: Compressor_14_3_F800_uid10
      port map ( X0 => Compressor_14_3_F800_uid10_bh3_uid163_In0,
                 X1 => Compressor_14_3_F800_uid10_bh3_uid163_In1,
                 R => Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164);
   Compressor_14_3_F800_uid10_bh3_uid163_Out0 <= Compressor_14_3_F800_uid10_bh3_uid163_Out0_copy164_d1; -- output copy to hold a pipeline register if needed

   bh3_w2_21 <= Compressor_14_3_F800_uid10_bh3_uid163_Out0(0);
   bh3_w3_18 <= Compressor_14_3_F800_uid10_bh3_uid163_Out0(1);
   bh3_w4_21 <= Compressor_14_3_F800_uid10_bh3_uid163_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid165_In0 <= "" & bh3_w4_20 & bh3_w4_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid165_In1 <= "" & bh3_w5_18 & bh3_w5_15;
   Compressor_23_3_F800_uid136_uid165: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid165_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid165_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166);
   Compressor_23_3_F800_uid136_bh3_uid165_Out0 <= Compressor_23_3_F800_uid136_bh3_uid165_Out0_copy166_d1; -- output copy to hold a pipeline register if needed

   bh3_w4_22 <= Compressor_23_3_F800_uid136_bh3_uid165_Out0(0);
   bh3_w5_19 <= Compressor_23_3_F800_uid136_bh3_uid165_Out0(1);
   bh3_w6_21 <= Compressor_23_3_F800_uid136_bh3_uid165_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid167_In0 <= "" & bh3_w6_20 & bh3_w6_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid167_In1 <= "" & bh3_w7_18 & bh3_w7_15;
   Compressor_23_3_F800_uid136_uid167: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid167_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid167_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168);
   Compressor_23_3_F800_uid136_bh3_uid167_Out0 <= Compressor_23_3_F800_uid136_bh3_uid167_Out0_copy168_d1; -- output copy to hold a pipeline register if needed

   bh3_w6_22 <= Compressor_23_3_F800_uid136_bh3_uid167_Out0(0);
   bh3_w7_19 <= Compressor_23_3_F800_uid136_bh3_uid167_Out0(1);
   bh3_w8_21 <= Compressor_23_3_F800_uid136_bh3_uid167_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid169_In0 <= "" & bh3_w8_20 & bh3_w8_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid169_In1 <= "" & bh3_w9_18 & bh3_w9_15;
   Compressor_23_3_F800_uid136_uid169: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid169_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid169_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170);
   Compressor_23_3_F800_uid136_bh3_uid169_Out0 <= Compressor_23_3_F800_uid136_bh3_uid169_Out0_copy170_d1; -- output copy to hold a pipeline register if needed

   bh3_w8_22 <= Compressor_23_3_F800_uid136_bh3_uid169_Out0(0);
   bh3_w9_19 <= Compressor_23_3_F800_uid136_bh3_uid169_Out0(1);
   bh3_w10_21 <= Compressor_23_3_F800_uid136_bh3_uid169_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid171_In0 <= "" & bh3_w10_20 & bh3_w10_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid171_In1 <= "" & bh3_w11_18 & bh3_w11_15;
   Compressor_23_3_F800_uid136_uid171: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid171_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid171_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172);
   Compressor_23_3_F800_uid136_bh3_uid171_Out0 <= Compressor_23_3_F800_uid136_bh3_uid171_Out0_copy172_d1; -- output copy to hold a pipeline register if needed

   bh3_w10_22 <= Compressor_23_3_F800_uid136_bh3_uid171_Out0(0);
   bh3_w11_19 <= Compressor_23_3_F800_uid136_bh3_uid171_Out0(1);
   bh3_w12_21 <= Compressor_23_3_F800_uid136_bh3_uid171_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid173_In0 <= "" & bh3_w12_20 & bh3_w12_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid173_In1 <= "" & bh3_w13_18 & bh3_w13_15;
   Compressor_23_3_F800_uid136_uid173: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid173_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid173_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174);
   Compressor_23_3_F800_uid136_bh3_uid173_Out0 <= Compressor_23_3_F800_uid136_bh3_uid173_Out0_copy174_d1; -- output copy to hold a pipeline register if needed

   bh3_w12_22 <= Compressor_23_3_F800_uid136_bh3_uid173_Out0(0);
   bh3_w13_19 <= Compressor_23_3_F800_uid136_bh3_uid173_Out0(1);
   bh3_w14_21 <= Compressor_23_3_F800_uid136_bh3_uid173_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid175_In0 <= "" & bh3_w14_20 & bh3_w14_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid175_In1 <= "" & bh3_w15_18 & bh3_w15_15;
   Compressor_23_3_F800_uid136_uid175: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid175_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid175_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176);
   Compressor_23_3_F800_uid136_bh3_uid175_Out0 <= Compressor_23_3_F800_uid136_bh3_uid175_Out0_copy176_d1; -- output copy to hold a pipeline register if needed

   bh3_w14_22 <= Compressor_23_3_F800_uid136_bh3_uid175_Out0(0);
   bh3_w15_19 <= Compressor_23_3_F800_uid136_bh3_uid175_Out0(1);
   bh3_w16_21 <= Compressor_23_3_F800_uid136_bh3_uid175_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid177_In0 <= "" & bh3_w16_20 & bh3_w16_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid177_In1 <= "" & bh3_w17_18 & bh3_w17_15;
   Compressor_23_3_F800_uid136_uid177: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid177_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid177_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178);
   Compressor_23_3_F800_uid136_bh3_uid177_Out0 <= Compressor_23_3_F800_uid136_bh3_uid177_Out0_copy178_d1; -- output copy to hold a pipeline register if needed

   bh3_w16_22 <= Compressor_23_3_F800_uid136_bh3_uid177_Out0(0);
   bh3_w17_19 <= Compressor_23_3_F800_uid136_bh3_uid177_Out0(1);
   bh3_w18_21 <= Compressor_23_3_F800_uid136_bh3_uid177_Out0(2);

   Compressor_23_3_F800_uid136_bh3_uid179_In0 <= "" & bh3_w18_20 & bh3_w18_19 & "0";
   Compressor_23_3_F800_uid136_bh3_uid179_In1 <= "" & bh3_w19_19 & bh3_w19_18;
   Compressor_23_3_F800_uid136_uid179: Compressor_23_3_F800_uid136
      port map ( X0 => Compressor_23_3_F800_uid136_bh3_uid179_In0,
                 X1 => Compressor_23_3_F800_uid136_bh3_uid179_In1,
                 R => Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180);
   Compressor_23_3_F800_uid136_bh3_uid179_Out0 <= Compressor_23_3_F800_uid136_bh3_uid179_Out0_copy180_d1; -- output copy to hold a pipeline register if needed

   bh3_w18_22 <= Compressor_23_3_F800_uid136_bh3_uid179_Out0(0);
   bh3_w19_20 <= Compressor_23_3_F800_uid136_bh3_uid179_Out0(1);
   bh3_w20_9 <= Compressor_23_3_F800_uid136_bh3_uid179_Out0(2);

   Compressor_3_2_F800_uid16_bh3_uid181_In0 <= "" & bh3_w20_8 & bh3_w20_7 & "0";
   Compressor_3_2_F800_uid16_uid181: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid181_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182);
   Compressor_3_2_F800_uid16_bh3_uid181_Out0 <= Compressor_3_2_F800_uid16_bh3_uid181_Out0_copy182_d1; -- output copy to hold a pipeline register if needed

   bh3_w20_10 <= Compressor_3_2_F800_uid16_bh3_uid181_Out0(0);
   bh3_w21_6 <= Compressor_3_2_F800_uid16_bh3_uid181_Out0(1);

   Compressor_3_2_F800_uid16_bh3_uid183_In0 <= "" & bh3_w21_5 & bh3_w21_4 & bh3_w21_3;
   Compressor_3_2_F800_uid16_uid183: Compressor_3_2_F800_uid16
      port map ( X0 => Compressor_3_2_F800_uid16_bh3_uid183_In0,
                 R => Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184);
   Compressor_3_2_F800_uid16_bh3_uid183_Out0 <= Compressor_3_2_F800_uid16_bh3_uid183_Out0_copy184_d1; -- output copy to hold a pipeline register if needed

   bh3_w21_7 <= Compressor_3_2_F800_uid16_bh3_uid183_Out0(0);
   bh3_w22_1 <= Compressor_3_2_F800_uid16_bh3_uid183_Out0(1);
   tmp_bitheapResult_bh3_3 <= bh3_w3_18 & bh3_w2_21 & bh3_w1_16_d1 & bh3_w0_13_d1;

   bitheapFinalAdd_bh3_In0 <= "0" & "0" & bh3_w22_0_d1 & bh3_w21_7 & bh3_w20_10 & bh3_w19_20 & bh3_w18_22 & bh3_w17_19 & bh3_w16_22 & bh3_w15_19 & bh3_w14_22 & bh3_w13_19 & bh3_w12_22 & bh3_w11_19 & bh3_w10_22 & bh3_w9_19 & bh3_w8_22 & bh3_w7_19 & bh3_w6_22 & bh3_w5_19 & bh3_w4_22;
   bitheapFinalAdd_bh3_In1 <= "0" & "0" & bh3_w22_1 & bh3_w21_6 & bh3_w20_9 & "0" & bh3_w18_21 & "0" & bh3_w16_21 & "0" & bh3_w14_21 & "0" & bh3_w12_21 & "0" & bh3_w10_21 & "0" & bh3_w8_21 & "0" & bh3_w6_21 & "0" & bh3_w4_21;
   bitheapFinalAdd_bh3_Cin <= '0';

   bitheapFinalAdd_bh3: IntAdder_21_F800_uid186
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh3_Cin,
                 X => bitheapFinalAdd_bh3_In0,
                 Y => bitheapFinalAdd_bh3_In1,
                 R => bitheapFinalAdd_bh3_Out);
   bitheapResult_bh3 <= bitheapFinalAdd_bh3_Out(19 downto 0) & tmp_bitheapResult_bh3_3_d2;
   OutRes <= bitheapResult_bh3;
   R <= OutRes;
end architecture;

